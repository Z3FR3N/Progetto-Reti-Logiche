//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "Prog_reti.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] in1;    //: /sn:0 {0}(#:-119,-555)(-119,-511){1}
//: {2}(-117,-509)(#:-86,-509){3}
//: {4}(-119,-507)(-119,-469)(-150,-469)(-150,-431){5}
reg [15:0] in3;    //: /sn:0 {0}(#:-300,-127)(-278,-127)(-278,-127)(-257,-127){1}
//: {2}(-255,-129)(-255,-168)(-401,-168)(#:-401,-555){3}
//: {4}(#:-255,-125)(#:-255,-85){5}
reg [7:0] in2;    //: /sn:0 {0}(#:-278,-509)(-245,-509){1}
//: {2}(-243,-511)(#:-243,-555){3}
//: {4}(-243,-507)(-243,-471)(-212,-471)(-212,-431){5}
wire [15:0] w13;    //: /sn:0 {0}(#:-216,34)(#:-216,6){1}
wire [15:0] w3;    //: /sn:0 {0}(#:-268,-311)(-217,-311){1}
//: {2}(-215,-313)(-215,-355){3}
//: {4}(-215,-309)(#:-215,-262){5}
wire [15:0] w12;    //: /sn:0 {0}(#:-298,-40)(#:-274,-40){1}
wire w10;    //: /sn:0 {0}(-255,-234)(-255,-220)(-230,-220){1}
wire [15:0] w1;    //: /sn:0 {0}(#:-150,-262)(-150,-309){1}
//: {2}(-148,-311)(-122,-311)(-122,-311)(#:-97,-311){3}
//: {4}(-150,-313)(-150,-355){5}
wire [15:0] w11;    //: /sn:0 {0}(#:-183,-85)(-183,-125){1}
//: {2}(-181,-127)(-170,-127)(-170,-127)(-164,-127){3}
//: {4}(-183,-129)(#:-183,-169){5}
//: enddecls

  //: LED g4 (w13) @(-216,41) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: joint g8 (in3) @(-255, -127) /w:[ -1 2 1 4 ]
  //: DIP g16 (in1) @(-119,-565) /sn:0 /w:[ 0 ] /st:128 /dn:1
  FD16 g3 (.B(in3), .A(w11), .R(w12), .Q(w13));   //: @(-273, -84) /sz:(109, 89) /R:3 /sn:0 /p:[ Ti0>5 Ti1>0 Lo0<1 Bo0<1 ]
  //: joint g17 (in1) @(-119, -509) /w:[ 2 1 -1 4 ]
  //: comment g26 @(-129,-218) /sn:0
  //: /line:"[A^2] + [B^2]"
  //: /end
  //: LED g2 (w3) @(-275,-311) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: comment g30 @(-157,47) /sn:0
  //: /line:"Q"
  //: /end
  //: joint g23 (w11) @(-183, -127) /w:[ 2 4 -1 1 ]
  RCA16 g1 (.B(w3), .A(w1), .Cout(w10), .S(w11));   //: @(-229, -261) /sz:(92, 91) /sn:0 /p:[ Ti0>5 Ti1>0 Lo0<1 Bo0<5 ]
  //: comment g24 @(-53,-340) /sn:0
  //: /line:"B^2"
  //: /end
  //: comment g29 @(-353,-156) /sn:0
  //: /line:"C"
  //: /end
  //: comment g18 @(-112,-156) /sn:0
  //: /line:"S"
  //: /end
  //: joint g10 (in2) @(-243, -509) /w:[ -1 2 1 4 ]
  //: comment g25 @(-332,-340) /sn:0
  //: /line:"A^2"
  //: /end
  //: DIP g6 (in3) @(-401,-565) /sn:0 /w:[ 3 ] /st:0 /dn:1
  //: joint g9 (w3) @(-215, -311) /w:[ -1 2 1 4 ]
  //: LED g7 (in3) @(-307,-127) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: comment g31 @(-412,-40) /sn:0
  //: /line:"R"
  //: /end
  //: LED g22 (w11) @(-157,-127) /sn:0 /R:3 /w:[ 3 ] /type:3
  //: DIP g12 (in2) @(-243,-565) /sn:0 /w:[ 3 ] /st:6 /dn:1
  //: comment g28 @(-313,-538) /sn:0
  //: /line:"A"
  //: /end
  POT2 g14 (.F(in1), .P(w1));   //: @(-175, -430) /sz:(53, 74) /sn:0 /p:[ Ti0>5 Bo0<5 ]
  //: LED g11 (w10) @(-255,-241) /sn:0 /w:[ 0 ] /type:0
  //: LED g5 (w12) @(-305,-40) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: comment g21 @(-57,-538) /sn:0
  //: /line:"B"
  //: /end
  //: LED g19 (in1) @(-79,-509) /sn:0 /R:3 /w:[ 3 ] /type:3
  //: LED g20 (w1) @(-90,-311) /sn:0 /R:3 /w:[ 3 ] /type:3
  //: joint g15 (w1) @(-150, -311) /w:[ 2 4 -1 1 ]
  POT2 g0 (.F(in2), .P(w3));   //: @(-241, -430) /sz:(56, 74) /sn:0 /p:[ Ti0>5 Bo0<3 ]
  //: comment g27 @(-153,-40) /sn:0
  //: /line:"{[A^2] + [B^2]} / C"
  //: /end
  //: LED g13 (in2) @(-285,-509) /sn:0 /R:1 /w:[ 0 ] /type:3

endmodule
//: /netlistEnd

//: /netlistBegin MUL16
module MUL16(B, P, A);
//: interface  /sz:(109, 40) /bd:[ Ti0>B[7:0](82/109) Ti1>A[7:0](18/109) Bo0<P[15:0](55/109) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] A;    //: /sn:0 {0}(#:857,243)(857,225){1}
//: {2}(857,224)(857,204){3}
//: {4}(857,203)(857,189){5}
//: {6}(857,188)(857,171){7}
//: {8}(857,170)(857,149){9}
//: {10}(857,148)(857,132){11}
//: {12}(857,131)(857,111){13}
//: {14}(857,110)(857,88){15}
//: {16}(#:857,87)(857,60){17}
input [7:0] B;    //: /sn:0 {0}(#:856,449)(856,423){1}
//: {2}(856,422)(856,402){3}
//: {4}(856,401)(856,383){5}
//: {6}(856,382)(856,366){7}
//: {8}(856,365)(856,350){9}
//: {10}(856,349)(856,331){11}
//: {12}(856,330)(856,312){13}
//: {14}(856,311)(856,295){15}
//: {16}(856,294)(#:856,281){17}
output [15:0] P;    //: /sn:0 {0}(900,2449)(#:852,2449){1}
wire w207;    //: /sn:0 {0}(-415,1255)(-415,1265)(-505,1265)(-505,1294){1}
wire P4;    //: /sn:0 {0}(30,1368)(30,2414)(846,2414){1}
wire w16;    //: /sn:0 {0}(-1144,1653)(-1144,1847){1}
wire w58;    //: /sn:0 {0}(293,718)(293,745)(235,745)(235,780){1}
wire w275;    //: /sn:0 {0}(-1609,2154)(-1722,2154){1}
wire w50;    //: /sn:0 {0}(255,549)(356,549){1}
wire P15;    //: /sn:0 {0}(-2006,2408)(-2013,2408)(-2013,2524)(846,2524){1}
wire P8;    //: /sn:0 {0}(-718,2444)(-718,2454)(846,2454){1}
wire w203;    //: /sn:0 {0}(-682,1613)(-562,1613){1}
wire B5;    //: {0}(-1448,1689)(0:-1448,1674)(-1267,1674){1}
//: {2}(1:-1263,1674)(-1043,1674){3}
//: {4}(2:-1039,1674)(-822,1674){5}
//: {6}(2:-818,1674)(-610,1674){7}
//: {8}(1:-608,1672)(-608,1539)(-544,1539)(-544,1413)(-400,1413){9}
//: {10}(1:-396,1413)(-235,1413){11}
//: {12}(3:-231,1413)(-41,1413){13}
//: {14}(1:-37,1413)(774,1413)(774,383)(851,383){15}
//: {16}(-39,1415)(-39,1428){17}
//: {18}(-233,1415)(-233,1428){19}
//: {20}(-398,1415)(-398,1428){21}
//: {22}(-608,1676)(-608,1692){23}
//: {24}(-820,1676)(-820,1688){25}
//: {26}(-1041,1676)(-1041,1689){27}
//: {28}(-1265,1676)(-1265,1689){29}
wire w4;    //: /sn:0 {0}(-1347,1653)(-1347,1847){1}
wire w39;    //: /sn:0 {0}(-491,435)(-491,463)(-514,463)(-514,511){1}
wire P6;    //: /sn:0 {0}(-331,1921)(-331,2434)(846,2434){1}
wire A3;    //: {0}(14:-1061,2223)(-1061,2083)(-924,2083)(-924,1942)(-848,1942){1}
//: {2}(1:-846,1940)(-846,1835)(-761,1835)(-761,1682)(-640,1682){3}
//: {4}(6:-638,1680)(-638,1587)(-586,1587)(-586,1146)(-434,1146){5}
//: {6}(8:-432,1144)(-432,1023)(-378,1023)(-378,870)(-248,870){7}
//: {8}(1:-246,868)(-246,782)(-192,782)(-192,605)(-68,605){9}
//: {10}(1:-66,603)(-66,171)(-33,171){11}
//: {12}(-29,171)(235,171){13}
//: {14}(239,171)(852,171){15}
//: {16}(94:237,173)(237,340){17}
//: {18}(94:-31,173)(-31,340){19}
//: {20}(-66,607)(-66,627){21}
//: {22}(-246,872)(-246,891){23}
//: {24}(-432,1148)(-432,1160){25}
//: {26}(-638,1684)(-638,1692){27}
//: {28}(-846,1944)(-846,1959){29}
wire w56;    //: /sn:0 {0}(261,818)(363,818){1}
wire w123;    //: /sn:0 {0}(-684,1068)(-564,1068){1}
wire w202;    //: /sn:0 {0}(-327,1107)(-327,1294){1}
wire w303;    //: /sn:0 {0}(-956,2193)(-956,2370){1}
wire w177;    //: /sn:0 {0}(-327,1371)(-327,1576){1}
wire w223;    //: /sn:0 {0}(-326,1653)(-326,1847){1}
wire w128;    //: /sn:0 {0}(-151,857)(-151,1030){1}
wire w189;    //: /sn:0 {0}(137,1243)(137,1265)(50,1265)(50,1294){1}
wire w0;    //: /sn:0 {0}(533,435)(533,476)(556,476)(556,511){1}
wire w132;    //: /sn:0 {0}(-506,2116)(-506,2061)(-424,2061)(-424,2054){1}
wire w22;    //: /sn:0 {0}(23,588)(23,780){1}
wire w20;    //: /sn:0 {0}(-708,1847)(-708,1799)(-625,1799)(-625,1787){1}
wire w261;    //: /sn:0 {0}(-724,1924)(-724,2116){1}
wire w30;    //: /sn:0 {0}(63,435)(63,475)(39,475)(39,511){1}
wire w196;    //: /sn:0 {0}(-148,1107)(-148,1294){1}
wire w185;    //: /sn:0 {0}(-59,1238)(-59,1264)(-132,1264)(-132,1294){1}
wire w122;    //: /sn:0 {0}(-480,1068)(-369,1068){1}
wire w42;    //: /sn:0 {0}(-14,435)(-14,473)(11,473)(11,511){1}
wire w218;    //: /sn:0 {0}(-478,1614)(-368,1614){1}
wire A6;    //: {0}(14:-1680,2223)(-1680,2071)(-1510,2071)(-1510,1935)(-1470,1935){1}
//: {2}(1:-1468,1933)(-1468,1815)(-1332,1815)(-1332,1668)(-1297,1668){3}
//: {4}(1:-1295,1666)(-1295,1574)(-1205,1574)(-1205,1393)(-1078,1393){5}
//: {6}(-1076,1391)(-1076,1288)(-1001,1288)(-1001,1123)(-858,1123){7}
//: {8}(1:-856,1121)(-856,1009)(-771,1009)(-771,870)(-649,870){9}
//: {10}(1:-647,868)(-647,788)(-609,788)(-609,290)(-584,290){11}
//: {12}(-582,288)(-582,111)(-317,111){13}
//: {14}(-313,111)(852,111){15}
//: {16}(94:-315,113)(-315,340){17}
//: {18}(99:-582,292)(-582,340){19}
//: {20}(-647,872)(-647,890){21}
//: {22}(-856,1125)(-856,1137)(-855,1137)(-855,1143){23}
//: {24}(18:-1076,1395)(-1076,1428){25}
//: {26}(-1295,1670)(-1295,1689){27}
//: {28}(-1468,1937)(-1468,1959){29}
wire w329;    //: /sn:0 {0}(-1303,2407)(-1182,2407){1}
wire w18;    //: /sn:0 {0}(-939,1847)(-939,1796)(-833,1796)(-833,1783){1}
wire w19;    //: /sn:0 {0}(-520,1653)(-520,1847){1}
wire A2;    //: {0}(10:-904,2223)(-904,2121)(-787,2121)(-787,1942)(-645,1942){1}
//: {2}(1:-643,1940)(-643,1809)(-573,1809)(-573,1403)(-430,1403){3}
//: {4}(1:-428,1401)(-428,1276)(-363,1276)(-363,1121)(-247,1121){5}
//: {6}(-245,1119)(-245,1019)(-188,1019)(-188,870)(-64,870){7}
//: {8}(1:-62,868)(-62,768)(-9,768)(-9,603)(116,603){9}
//: {10}(1:118,601)(118,189)(157,189){11}
//: {12}(161,189)(418,189){13}
//: {14}(422,189)(852,189){15}
//: {16}(93:420,191)(420,340){17}
//: {18}(159,191)(7:159,340){19}
//: {20}(118,605)(118,627){21}
//: {22}(-62,872)(-62,891){23}
//: {24}(26:-245,1123)(-245,1149){25}
//: {26}(-428,1405)(-428,1428){27}
//: {28}(-643,1944)(-643,1966){29}
wire w12;    //: /sn:0 {0}(437,435)(437,475)(414,475)(414,511){1}
wire w190;    //: /sn:0 {0}(-1102,1614)(-991,1614){1}
wire B2;    //: {0}(-798,891)(1:-798,876)(-619,876){1}
//: {2}(1:-617,874)(-617,802)(-599,802)(-599,612)(-411,612){3}
//: {4}(1:-407,612)(-241,612){5}
//: {6}(3:-237,612)(-38,612){7}
//: {8}(1:-34,612)(146,612){9}
//: {10}(1:150,612)(308,612){11}
//: {12}(1:312,612)(510,612){13}
//: {14}(4:514,612)(730,612)(730,331)(851,331){15}
//: {16}(512,614)(512,627){17}
//: {18}(310,614)(310,623){19}
//: {20}(148,614)(148,627){21}
//: {22}(-36,614)(-36,627){23}
//: {24}(-239,614)(-239,629){25}
//: {26}(-409,614)(-409,628){27}
//: {28}(-617,878)(-617,890){29}
wire B7;    //: {0}(99:-1878,2223)(-1878,2211)(-1652,2211){1}
//: {2}(2:-1648,2211)(-1440,2211){3}
//: {4}(1:-1436,2211)(-1255,2211){5}
//: {6}(4:-1251,2211)(-1033,2211){7}
//: {8}(11:-1029,2211)(-876,2211){9}
//: {10}(1:-872,2211)(-616,2211){11}
//: {12}(5:-612,2211)(-571,2211)(-571,1942)(-413,1942){13}
//: {14}(0:-409,1942)(798,1942)(798,423)(851,423){15}
//: {16}(-411,1944)(-411,1959){17}
//: {18}(-614,2213)(-614,2223){19}
//: {20}(-874,2213)(-874,2223){21}
//: {22}(-1031,2213)(-1031,2223){23}
//: {24}(-1253,2213)(-1253,2223){25}
//: {26}(-1438,2213)(-1438,2223){27}
//: {28}(-1650,2213)(-1650,2223){29}
wire w54;    //: /sn:0 {0}(499,722)(499,743)(418,743)(418,780){1}
wire w269;    //: /sn:0 {0}(-708,1576)(-708,1538)(-631,1538)(-631,1524){1}
wire w335;    //: /sn:0 {0}(-1455,2318)(-1455,2333)(-1551,2333)(-1551,2370){1}
wire w180;    //: /sn:0 {0}(219,1032)(219,857){1}
wire w86;    //: /sn:0 {0}(-730,857)(-730,1030){1}
wire w31;    //: /sn:0 {0}(27,1032)(27,857){1}
wire w247;    //: /sn:0 {0}(-955,1924)(-955,2116){1}
wire B1;    //: {0}(5:-632,628)(-632,312)(-554,312){1}
//: {2}(-1:-550,312)(-357,312){3}
//: {4}(-353,312)(-180,312){5}
//: {6}(-176,312)(-3,312){7}
//: {8}(1,312)(187,312){9}
//: {10}(191,312)(375,312){11}
//: {12}(379,312)(544,312){13}
//: {14}(548,312)(851,312){15}
//: {16}(57:546,314)(546,340){17}
//: {18}(61:377,314)(377,340){19}
//: {20}(65:189,314)(189,340){21}
//: {22}(61:-1,314)(-1,340){23}
//: {24}(50:-178,314)(-178,340){25}
//: {26}(99:-355,314)(-355,340){27}
//: {28}(-552,314)(-552,340){29}
wire w199;    //: /sn:0 {0}(-228,1244)(-228,1261)(-311,1261)(-311,1294){1}
wire w116;    //: /sn:0 {0}(-106,1068)(-12,1068){1}
wire P14;    //: /sn:0 {0}(-1964,2447)(-1964,2514)(846,2514){1}
wire w110;    //: /sn:0 {0}(-772,818)(-949,818)(-949,1030){1}
wire w8;    //: /sn:0 {0}(-1461,1784)(-1461,1793)(-1542,1793)(-1542,1847){1}
wire w115;    //: /sn:0 {0}(72,1070)(186,1070){1}
wire w140;    //: /sn:0 {0}(-707,2116)(-707,2074)(-630,2074)(-630,2061){1}
wire w233;    //: /sn:0 {0}(-1390,1885)(-1518,1885){1}
wire P5;    //: /sn:0 {0}(-152,1650)(-152,2424)(846,2424){1}
wire B6;    //: {0}(-1641,1959)(0:-1641,1947)(-1440,1947){1}
//: {2}(1:-1436,1947)(-1257,1947){3}
//: {4}(6:-1253,1947)(-1039,1947){5}
//: {6}(1:-1035,1947)(-818,1947){7}
//: {8}(1:-814,1947)(-615,1947){9}
//: {10}(1:-613,1945)(-613,1822)(-565,1822)(-565,1676)(-409,1676){11}
//: {12}(2:-405,1676)(-227,1676){13}
//: {14}(0:-223,1676)(787,1676)(787,402)(851,402){15}
//: {16}(-225,1678)(-225,1691){17}
//: {18}(-407,1678)(-407,1689){19}
//: {20}(-613,1949)(-613,1966){21}
//: {22}(-816,1949)(-816,1959){23}
//: {24}(-1037,1949)(-1037,1959){25}
//: {26}(-1255,1949)(-1255,1959){27}
//: {28}(-1438,1949)(-1438,1959){29}
wire w276;    //: /sn:0 {0}(-1566,2193)(-1566,2370){1}
wire w260;    //: /sn:0 {0}(-682,1885)(-562,1885){1}
wire w136;    //: /sn:0 {0}(-285,1067)(-190,1067){1}
wire w35;    //: /sn:0 {0}(-530,588)(-530,780){1}
wire w67;    //: /sn:0 {0}(-1654,2054)(-1654,2065)(-1744,2065)(-1744,2116){1}
wire w28;    //: /sn:0 {0}(-313,1847)(-313,1796)(-242,1796)(-242,1786){1}
wire w169;    //: /sn:0 {0}(-726,1107)(-726,1294){1}
wire w135;    //: /sn:0 {0}(-430,991)(-430,997)(-506,997)(-506,1030){1}
wire w346;    //: /sn:0 {0}(-891,2318)(-891,2326)(-935,2326)(-935,2370){1}
wire w14;    //: /sn:0 {0}(-1127,1847)(-1127,1807)(-1058,1807)(-1058,1784){1}
wire w45;    //: /sn:0 {0}(-368,435)(-368,466)(-345,466)(-345,511){1}
wire w204;    //: /sn:0 {0}(-907,1614)(-766,1614){1}
wire w11;    //: /sn:0 {0}(-1282,1784)(-1282,1824)(-1332,1824)(-1332,1847){1}
wire w78;    //: /sn:0 {0}(-525,857)(-525,1030){1}
wire w74;    //: /sn:0 {0}(-483,818)(-372,818){1}
wire w2;    //: /sn:0 {0}(440,549)(537,549){1}
wire P13;    //: /sn:0 {0}(-1771,2447)(-1771,2504)(846,2504){1}
wire w274;    //: /sn:0 {0}(-1523,2151)(-1390,2151){1}
wire A7;    //: {0}(7:-1908,2223)(-1908,1931)(-1673,1931){1}
//: {2}(-1671,1929)(-1671,1640)(-1480,1640){3}
//: {4}(-1478,1638)(-1478,1389)(-1291,1389){5}
//: {6}(-1289,1387)(-1289,1100)(-1065,1100){7}
//: {8}(-1063,1098)(-1063,839)(-830,839){9}
//: {10}(-828,837)(-828,581)(-664,581){11}
//: {12}(-662,579)(-662,88)(-510,88){13}
//: {14}(-506,88)(852,88){15}
//: {16}(94:-508,90)(-508,340){17}
//: {18}(33:-662,583)(-662,628){19}
//: {20}(72:-828,841)(-828,891){21}
//: {22}(55:-1063,1102)(-1063,1149){23}
//: {24}(24:-1289,1391)(-1289,1428){25}
//: {26}(57:-1478,1642)(-1478,1689){27}
//: {28}(19:-1671,1933)(-1671,1959){29}
wire P10;    //: /sn:0 {0}(-1140,2447)(-1140,2474)(846,2474){1}
wire w105;    //: /sn:0 {0}(319,986)(319,997)(241,997)(241,1032){1}
wire A1;    //: {0}(15:-644,2223)(-644,2089)(-580,2089)(-580,1841)(-544,1841)(-544,1667)(-439,1667){1}
//: {2}(-437,1665)(-437,1578)(-371,1578)(-371,1399)(-265,1399){3}
//: {4}(-263,1397)(-263,1273)(-188,1273)(-188,1123)(-74,1123){5}
//: {6}(1:-72,1121)(-72,1012)(-10,1012)(-10,865)(110,865){7}
//: {8}(1:112,863)(112,769)(178,769)(178,602)(278,602){9}
//: {10}(280,600)(280,510)(305,510)(305,204)(345,204){11}
//: {12}(349,204)(592,204){13}
//: {14}(596,204)(852,204){15}
//: {16}(90:594,206)(594,340){17}
//: {18}(347,206)(8:347,340){19}
//: {20}(31:280,604)(280,623){21}
//: {22}(112,867)(112,887){23}
//: {24}(-72,1125)(-72,1143){25}
//: {26}(33:-263,1401)(-263,1428){27}
//: {28}(26:-437,1669)(-437,1689){29}
wire w228;    //: /sn:0 {0}(-478,1885)(-368,1885){1}
wire w288;    //: /sn:0 {0}(-1306,2154)(-1180,2154){1}
wire w15;    //: /sn:0 {0}(364,435)(364,474)(386,474)(386,511){1}
wire w55;    //: /sn:0 {0}(213,588)(213,780){1}
wire B4;    //: {0}(-1259,1428)(1:-1259,1411)(-1048,1411){1}
//: {2}(2:-1044,1411)(-829,1411){3}
//: {4}(2:-825,1411)(-616,1411){5}
//: {6}(1:-614,1409)(-614,1289)(-563,1289)(-563,1134)(-404,1134){7}
//: {8}(1:-400,1134)(-217,1134){9}
//: {10}(1:-213,1134)(-44,1134){11}
//: {12}(1:-40,1134)(148,1134){13}
//: {14}(1:152,1134)(761,1134)(761,366)(851,366){15}
//: {16}(150,1136)(150,1148){17}
//: {18}(-42,1136)(-42,1143){19}
//: {20}(-215,1136)(-215,1149){21}
//: {22}(-402,1136)(-402,1160){23}
//: {24}(-614,1413)(-614,1429){25}
//: {26}(-827,1413)(-827,1428){27}
//: {28}(-1046,1413)(-1046,1428){29}
wire w92;    //: /sn:0 {0}(-45,986)(-45,998)(-132,998)(-132,1030){1}
wire w94;    //: /sn:0 {0}(-979,1068)(-1155,1068)(-1155,1294){1}
wire w87;    //: /sn:0 {0}(125,982)(125,998)(46,998)(46,1032){1}
wire w76;    //: /sn:0 {0}(-426,723)(-426,746)(-504,746)(-504,780){1}
wire B0;    //: {0}(37:-478,340)(-478,295)(-287,295){1}
//: {2}(-283,295)(-106,295){3}
//: {4}(-102,295)(74,295){5}
//: {6}(78,295)(265,295){7}
//: {8}(269,295)(448,295){9}
//: {10}(452,295)(622,295){11}
//: {12}(626,295)(705,295){13}
//: {14}(709,295)(851,295){15}
//: {16}(76:707,297)(707,340){17}
//: {18}(74:624,297)(624,340){19}
//: {20}(81:450,297)(450,340){21}
//: {22}(81:267,297)(267,340){23}
//: {24}(74:76,297)(76,340){25}
//: {26}(79:-104,297)(-104,340){27}
//: {28}(74:-285,297)(-285,340){29}
wire w172;    //: /sn:0 {0}(-1185,1332)(-1359,1332)(-1359,1576){1}
wire w286;    //: /sn:0 {0}(-1050,2054)(-1050,2069)(-1122,2069)(-1122,2116){1}
wire w183;    //: /sn:0 {0}(30,1109)(30,1294){1}
wire w114;    //: /sn:0 {0}(-109,817)(-15,817){1}
wire w262;    //: /sn:0 {0}(-134,1576)(-134,1534)(-52,1534)(-52,1523){1}
wire A0;    //: {0}(12:-441,1959)(-441,1826)(-364,1826)(-364,1666)(-257,1666){1}
//: {2}(1:-255,1664)(-255,1562)(-192,1562)(-192,1401)(-71,1401){3}
//: {4}(1:-69,1399)(-69,1280)(2,1280)(2,1125)(116,1125){5}
//: {6}(118,1123)(118,1010)(178,1010)(178,870)(300,870){7}
//: {8}(1:302,868)(302,763)(355,763)(355,603)(480,603){9}
//: {10}(482,601)(482,225)(514,225){11}
//: {12}(518,225)(675,225){13}
//: {14}(679,225)(852,225){15}
//: {16}(92:677,227)(677,340){17}
//: {18}(92:516,227)(516,340){19}
//: {20}(18:482,605)(482,627){21}
//: {22}(302,872)(302,891){23}
//: {24}(28:118,1127)(118,1148){25}
//: {26}(-69,1403)(-69,1428){27}
//: {28}(-255,1668)(-255,1691){29}
wire w307;    //: /sn:0 {0}(-723,2193)(-723,2370){1}
wire w6;    //: /sn:0 {0}(-375,549)(-488,549){1}
wire w65;    //: /sn:0 {0}(-49,722)(-49,746)(-135,746)(-135,780){1}
wire w264;    //: /sn:0 {0}(-504,1576)(-504,1536)(-411,1536)(-411,1523){1}
wire w344;    //: /sn:0 {0}(-1098,2408)(-993,2408){1}
wire w291;    //: /sn:0 {0}(-1272,2054)(-1272,2082)(-1332,2082)(-1332,2116){1}
wire A5;    //: {0}(21:-1468,2223)(-1468,2136)(-1403,2136)(-1403,1937)(-1287,1937){1}
//: {2}(1:-1285,1935)(-1285,1868)(-1237,1868)(-1237,1667)(-1073,1667){3}
//: {4}(1:-1071,1665)(-1071,1560)(-1013,1560)(-1013,1394)(-859,1394){5}
//: {6}(-857,1392)(-857,1319)(-788,1319)(-788,1120)(-659,1120){7}
//: {8}(1:-657,1118)(-657,1009)(-591,1009)(-591,602)(-441,602){9}
//: {10}(1:-439,600)(-439,132)(-387,132){11}
//: {12}(-383,132)(-136,132){13}
//: {14}(-132,132)(852,132){15}
//: {16}(93:-134,134)(-134,340){17}
//: {18}(97:-385,134)(-385,340){19}
//: {20}(-439,604)(-439,628){21}
//: {22}(-657,1122)(-657,1151){23}
//: {24}(37:-857,1396)(-857,1428){25}
//: {26}(-1071,1669)(-1071,1689){27}
//: {28}(-1285,1939)(-1285,1959){29}
wire w59;    //: /sn:0 {0}(-291,549)(-243,549)(-243,549)(-200,549){1}
wire w205;    //: /sn:0 {0}(-724,1653)(-724,1847){1}
wire w252;    //: /sn:0 {0}(-1143,1924)(-1143,2116){1}
wire w25;    //: /sn:0 {0}(-504,1847)(-504,1800)(-414,1800)(-414,1784){1}
wire P1;    //: /sn:0 {0}(574,585)(574,2384)(846,2384){1}
wire w62;    //: /sn:0 {0}(254,435)(254,472)(229,472)(229,511){1}
wire w306;    //: /sn:0 {0}(-1667,2318)(-1667,2333)(-1755,2333)(-1755,2370){1}
wire w337;    //: /sn:0 {0}(-1044,2318)(-1044,2329)(-1124,2329)(-1124,2370){1}
wire w241;    //: /sn:0 {0}(-725,1371)(-725,1576){1}
wire w162;    //: /sn:0 {0}(-683,1332)(-563,1332){1}
wire w186;    //: /sn:0 {0}(-284,1614)(-189,1614){1}
wire w159;    //: /sn:0 {0}(-1046,1244)(-1046,1251)(-1123,1251)(-1123,1294){1}
wire w176;    //: /sn:0 {0}(-285,1332)(-190,1332){1}
wire w142;    //: /sn:0 {0}(-634,985)(-634,997)(-710,997)(-710,1030){1}
wire w299;    //: /sn:0 {0}(-1764,2193)(-1764,2370){1}
wire w36;    //: /sn:0 {0}(-191,435)(-191,474)(-170,474)(-170,511){1}
wire w82;    //: /sn:0 {0}(-645,723)(-645,748)(-714,748)(-714,780){1}
wire w60;    //: /sn:0 {0}(69,818)(177,818){1}
wire w225;    //: /sn:0 {0}(-1128,1576)(-1128,1536)(-1063,1536)(-1063,1523){1}
wire w124;    //: /sn:0 {0}(-522,1107)(-522,1294){1}
wire w148;    //: /sn:0 {0}(-900,1332)(-767,1332){1}
wire w112;    //: /sn:0 {0}(-842,1238)(-842,1255)(-926,1255)(-926,1294){1}
wire w234;    //: /sn:0 {0}(-1348,1924)(-1348,2116){1}
wire w37;    //: /sn:0 {0}(-333,588)(-333,780){1}
wire w255;    //: /sn:0 {0}(-148,1371)(-148,1576){1}
wire w214;    //: /sn:0 {0}(-1389,1614)(-1576,1614)(-1576,1847){1}
wire w73;    //: /sn:0 {0}(-256,724)(-256,758)(-314,758)(-314,780){1}
wire w217;    //: /sn:0 {0}(-1327,1576)(-1327,1538)(-1272,1538)(-1272,1523){1}
wire w211;    //: /sn:0 {0}(-709,1294)(-709,1257)(-644,1257)(-644,1246){1}
wire w63;    //: /sn:0 {0}(-949,1653)(-949,1847){1}
wire w270;    //: /sn:0 {0}(-681,2154)(-561,2154){1}
wire w70;    //: /sn:0 {0}(135,722)(135,745)(43,745)(43,780){1}
wire w111;    //: /sn:0 {0}(-768,1068)(-895,1068){1}
wire w21;    //: /sn:0 {0}(176,435)(176,473)(201,473)(201,511){1}
wire w24;    //: /sn:0 {0}(-298,435)(-298,465)(-317,465)(-317,511){1}
wire w256;    //: /sn:0 {0}(-1607,1885)(-1776,1885)(-1776,2116){1}
wire w302;    //: /sn:0 {0}(-914,2154)(-765,2154){1}
wire w246;    //: /sn:0 {0}(-1101,1885)(-997,1885){1}
wire w287;    //: /sn:0 {0}(-1096,2153)(-998,2153){1}
wire w317;    //: /sn:0 {0}(-1813,2408)(-1922,2408){1}
wire w304;    //: /sn:0 {0}(-1891,2318)(-1891,2330)(-1944,2330)(-1944,2370){1}
wire w224;    //: /sn:0 {0}(-310,1576)(-310,1540)(-250,1540)(-250,1523){1}
wire P3;    //: /sn:0 {0}(223,1106)(223,2404)(846,2404){1}
wire w144;    //: /sn:0 {0}(-917,1030)(-917,996)(-811,996)(-811,986){1}
wire w316;    //: /sn:0 {0}(-1729,2408)(-1609,2408){1}
wire w52;    //: /sn:0 {0}(65,548)(171,548){1}
wire w232;    //: /sn:0 {0}(-1306,1885)(-1185,1885){1}
wire w191;    //: /sn:0 {0}(-1186,1614)(-1305,1614){1}
wire w75;    //: /sn:0 {0}(-567,818)(-688,818){1}
wire w150;    //: /sn:0 {0}(-942,1371)(-942,1576){1}
wire P7;    //: /sn:0 {0}(-524,2190)(-524,2444)(846,2444){1}
wire w17;    //: /sn:0 {0}(-158,588)(-158,780){1}
wire w330;    //: /sn:0 {0}(-1525,2408)(-1387,2408){1}
wire w33;    //: /sn:0 {0}(-117,435)(-117,476)(-142,476)(-142,511){1}
wire P12;    //: /sn:0 {0}(-1567,2447)(-1567,2494)(846,2494){1}
wire w145;    //: /sn:0 {0}(-106,1332)(-11,1332){1}
wire w49;    //: /sn:0 {0}(611,435)(611,475)(592,475)(592,511){1}
wire P11;    //: /sn:0 {0}(-1345,2447)(-1345,2484)(846,2484){1}
wire w48;    //: /sn:0 {0}(-565,435)(-565,463)(-542,463)(-542,511){1}
wire w257;    //: /sn:0 {0}(-1563,1924)(-1563,2116){1}
wire w47;    //: /sn:0 {0}(398,588)(398,780){1}
wire w294;    //: /sn:0 {0}(-1348,2193)(-1348,2370){1}
wire w149;    //: /sn:0 {0}(-984,1332)(-1101,1332){1}
wire w280;    //: /sn:0 {0}(-829,2054)(-829,2097)(-940,2097)(-940,2116){1}
wire w245;    //: /sn:0 {0}(-913,1884)(-766,1884){1}
wire w161;    //: /sn:0 {0}(-479,1331)(-369,1331){1}
wire w85;    //: /sn:0 {0}(-229,986)(-229,999)(-311,999)(-311,1030){1}
wire w90;    //: /sn:0 {0}(-288,818)(-193,818){1}
wire w289;    //: /sn:0 {0}(-1138,2193)(-1138,2370){1}
wire w267;    //: /sn:0 {0}(-521,1371)(-521,1576){1}
wire B3;    //: {0}(-1033,1149)(0:-1033,1130)(-827,1130){1}
//: {2}(3:-823,1130)(-629,1130){3}
//: {4}(1:-627,1128)(-627,1017)(-583,1017)(-583,876)(-415,876){5}
//: {6}(3:-411,876)(-218,876){7}
//: {8}(3:-214,876)(-34,876){9}
//: {10}(3:-30,876)(140,876){11}
//: {12}(4:144,876)(330,876){13}
//: {14}(1:334,876)(745,876)(745,350)(851,350){15}
//: {16}(332,878)(332,891){17}
//: {18}(142,878)(142,887){19}
//: {20}(-32,878)(-32,891){21}
//: {22}(-216,878)(-216,891){23}
//: {24}(-413,878)(-413,896){25}
//: {26}(-627,1132)(-627,1151){27}
//: {28}(-825,1132)(-825,1143){29}
wire P0;    //: /sn:0 {0}(694,435)(694,2374)(846,2374){1}
wire w5;    //: /sn:0 {0}(-1266,2318)(-1266,2326)(-1329,2326)(-1329,2370){1}
wire w350;    //: /sn:0 {0}(-627,2318)(-627,2341)(-700,2341)(-700,2370){1}
wire w9;    //: /sn:0 {0}(-116,549)(-19,549){1}
wire w265;    //: /sn:0 {0}(-520,1924)(-520,2116){1}
wire A4;    //: {0}(15:-1283,2223)(-1283,2101)(-1213,2101)(-1213,1938)(-1069,1938){1}
//: {2}(1:-1067,1936)(-1067,1848)(-1010,1848)(-1010,1667)(-852,1667){3}
//: {4}(1:-850,1665)(-850,1567)(-781,1567)(-781,1403)(-646,1403){5}
//: {6}(1:-644,1401)(-644,1277)(-575,1277)(-575,884)(-445,884){7}
//: {8}(8:-443,882)(-443,771)(-373,771)(-373,602)(-271,602){9}
//: {10}(1:-269,600)(-269,521)(-249,521)(-249,149)(-210,149){11}
//: {12}(-206,149)(44,149){13}
//: {14}(48,149)(852,149){15}
//: {16}(93:46,151)(46,340){17}
//: {18}(-208,151)(6:-208,340){19}
//: {20}(-269,604)(-269,629){21}
//: {22}(-443,886)(-443,896){23}
//: {24}(-644,1405)(-644,1429){25}
//: {26}(-850,1669)(-850,1688){27}
//: {28}(-1067,1940)(-1067,1959){29}
wire w220;    //: /sn:0 {0}(-1143,1371)(-1143,1576){1}
wire w231;    //: /sn:0 {0}(-933,1576)(-933,1547)(-844,1547)(-844,1523){1}
wire P2;    //: /sn:0 {0}(400,854)(400,2394)(846,2394){1}
wire w312;    //: /sn:0 {0}(-909,2408)(-755,2408){1}
wire w298;    //: /sn:0 {0}(-1806,2154)(-1976,2154)(-1976,2191)(-1976,2191)(-1976,2370){1}
wire w301;    //: /sn:0 {0}(-1455,2054)(-1455,2095)(-1550,2095)(-1550,2116){1}
wire w157;    //: /sn:0 {0}(-937,1107)(-937,1294){1}
wire w93;    //: /sn:0 {0}(-330,857)(-330,1030){1}
wire P9;    //: /sn:0 {0}(-951,2447)(-951,2464)(846,2464){1}
wire w77;    //: /sn:0 {0}(-572,549)(-742,549)(-742,780){1}
//: enddecls

  //: joint g246 (A4) @(-1067, 1938) /w:[ -1 2 1 28 ]
  //: joint g164 (B3) @(332, 876) /w:[ 14 -1 13 16 ]
  NandAND g8 (.in2(A2), .in1(B0), .out(w12));   //: @(400, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>21 Bo0<0 ]
  FA g4 (.b(w12), .a(w15), .Cin(w2), .Cout(w50), .S(w47));   //: @(357, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g116 (.b(w335), .a(w276), .Cin(w330), .Cout(w316), .S(P12));   //: @(-1608, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g197 (A0) @(118, 1125) /w:[ -1 6 5 24 ]
  assign A0 = A[0]; //: TAP g157 @(855,225) /sn:0 /R:2 /w:[ 15 1 2 ] /ss:0
  //: joint g224 (B6) @(-407, 1676) /w:[ 12 -1 11 18 ]
  NandAND g17 (.in2(A5), .in1(B0), .out(w33));   //: @(-154, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>27 Bo0<0 ]
  //: joint g243 (A1) @(-437, 1667) /w:[ -1 2 1 28 ]
  //: joint g226 (B6) @(-816, 1947) /w:[ 8 -1 7 22 ]
  //: joint g137 (B0) @(-104, 295) /w:[ 4 -1 3 26 ]
  //: joint g198 (A1) @(-72, 1123) /w:[ -1 6 5 24 ]
  NandAND g92 (.in2(B5), .in1(A6), .out(w11));   //: @(-1309, 1690) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>27 Bo0<0 ]
  NandAND g30 (.in2(B2), .in1(A4), .out(w73));   //: @(-283, 630) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>21 Bo0<0 ]
  FA g74 (.b(w231), .a(w150), .Cin(w204), .Cout(w190), .S(w63));   //: @(-990, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g130 (B1) @(377, 312) /w:[ 12 -1 11 18 ]
  assign A5 = A[5]; //: TAP g183 @(855,132) /sn:0 /R:2 /w:[ 15 11 12 ] /ss:0
  //: IN g1 (B) @(856,279) /sn:0 /R:3 /w:[ 17 ]
  FA g77 (.b(w264), .a(w267), .Cin(w218), .Cout(w203), .S(w19));   //: @(-561, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g214 (B5) @(-820, 1674) /w:[ 6 -1 5 24 ]
  NandAND g111 (.in2(A3), .in1(B7), .out(w337));   //: @(-1081, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>23 Bo0<0 ]
  //: joint g179 (B4) @(-215, 1134) /w:[ 10 -1 9 20 ]
  //: joint g144 (B2) @(148, 612) /w:[ 10 -1 9 20 ]
  NandAND g51 (.in2(B3), .in1(A1), .out(w87));   //: @(98, 888) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>23 Bo0<0 ]
  //: joint g206 (A6) @(-856, 1123) /w:[ -1 8 7 22 ]
  //: joint g190 (B3) @(-825, 1130) /w:[ 2 -1 1 28 ]
  //: joint g161 (B3) @(142, 876) /w:[ 12 -1 11 18 ]
  NandAND g70 (.in2(B4), .in1(A5), .out(w231));   //: @(-871, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>25 Bo0<1 ]
  //: joint g149 (A2) @(159, 189) /w:[ 12 -1 11 18 ]
  NandAND g103 (.in2(A4), .in1(B6), .out(w286));   //: @(-1087, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>25 Bo0<0 ]
  NandAND g25 (.in2(A0), .in1(B2), .out(w54));   //: @(462, 628) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>17 Bo0<0 ]
  NandAND g10 (.in2(A1), .in1(B1), .out(w15));   //: @(327, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>19 Bo0<0 ]
  FA g65 (.b(w185), .a(w196), .Cin(w145), .Cout(w176), .S(w255));   //: @(-189, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g220 (A6) @(-1076, 1393) /w:[ -1 6 5 24 ]
  NandAND g64 (.in2(B3), .in1(A6), .out(w112));   //: @(-869, 1144) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>23 Bo0<0 ]
  //: joint g185 (A1) @(112, 865) /w:[ -1 8 7 22 ]
  NandAND g49 (.in2(B2), .in1(A6), .out(w142));   //: @(-661, 891) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>21 Bo0<0 ]
  FA g72 (.b(w269), .a(w241), .Cin(w203), .Cout(w204), .S(w205));   //: @(-765, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: OUT g251 (P) @(897,2449) /sn:0 /w:[ 0 ]
  //: joint g142 (B1) @(-355, 312) /w:[ 4 -1 3 26 ]
  //: joint g136 (B1) @(-1, 312) /w:[ 8 -1 7 22 ]
  NandAND g6 (.in2(A1), .in1(B0), .out(w49));   //: @(574, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>19 Bo0<0 ]
  assign B1 = B[1]; //: TAP g124 @(854,312) /sn:0 /R:2 /w:[ 15 13 14 ] /ss:0
  NandAND g56 (.in2(B3), .in1(A5), .out(w211));   //: @(-671, 1152) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>23 Bo0<1 ]
  NandAND g7 (.in2(A0), .in1(B1), .out(w0));   //: @(496, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>17 Bo0<0 ]
  FA g35 (.b(w82), .a(w77), .Cin(w75), .Cout(w110), .S(w86));   //: @(-771, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g58 (.b(w207), .a(w124), .Cin(w161), .Cout(w162), .S(w267));   //: @(-562, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g229 (B6) @(-1438, 1947) /w:[ 2 -1 1 28 ]
  //: joint g200 (B4) @(-402, 1134) /w:[ 8 -1 7 22 ]
  NandAND g98 (.in2(B6), .in1(A5), .out(w291));   //: @(-1299, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>29 Bo0<0 ]
  assign A4 = A[4]; //: TAP g181 @(855,149) /sn:0 /R:2 /w:[ 15 9 10 ] /ss:0
  //: joint g204 (A7) @(-1063, 1100) /w:[ -1 8 7 22 ]
  //: joint g192 (A6) @(-647, 870) /w:[ -1 10 9 20 ]
  NandAND g85 (.in2(A7), .in1(B5), .out(w8));   //: @(-1498, 1690) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  HA g67 (.b(w262), .a(w255), .Cout(w186), .S(P5));   //: @(-188, 1577) /sz:(72, 72) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<1 Bo0<0 ]
  //: joint g126 (B1) @(546, 312) /w:[ 14 -1 13 16 ]
  //: joint g234 (A6) @(-1295, 1668) /w:[ -1 4 3 26 ]
  //: joint g208 (B6) @(-225, 1676) /w:[ 14 -1 13 16 ]
  HA g33 (.b(w54), .a(w47), .Cout(w56), .S(P2));   //: @(364, 781) /sz:(72, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  FA g54 (.b(w112), .a(w157), .Cin(w148), .Cout(w149), .S(w150));   //: @(-983, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  NandAND g40 (.in2(B3), .in1(A4), .out(w135));   //: @(-457, 897) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>23 Bo0<0 ]
  FA g52 (.b(w92), .a(w128), .Cin(w116), .Cout(w136), .S(w196));   //: @(-189, 1031) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  HA g81 (.b(w28), .a(w223), .Cout(w228), .S(P6));   //: @(-367, 1848) /sz:(72, 72) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<1 Bo0<0 ]
  //: joint g163 (B3) @(-216, 876) /w:[ 8 -1 7 22 ]
  //: joint g132 (A3) @(237, 171) /w:[ 14 -1 13 16 ]
  assign B7 = B[7]; //: TAP g222 @(854,423) /sn:0 /R:2 /w:[ 15 1 2 ] /ss:0
  //: joint g217 (A3) @(-432, 1146) /w:[ -1 6 5 24 ]
  //: joint g210 (A0) @(-69, 1401) /w:[ -1 4 3 26 ]
  NandAND g108 (.in2(B6), .in1(A2), .out(w140));   //: @(-657, 1967) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>29 Bo0<1 ]
  NandAND g12 (.in2(A2), .in1(B1), .out(w21));   //: @(139, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>21 Bo0<0 ]
  //: joint g131 (B0) @(267, 295) /w:[ 8 -1 7 22 ]
  NandAND g106 (.in2(B6), .in1(A6), .out(w301));   //: @(-1482, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>29 Bo0<0 ]
  //: joint g230 (A2) @(-428, 1403) /w:[ -1 4 3 26 ]
  //: joint g194 (B5) @(-233, 1413) /w:[ 12 -1 11 18 ]
  //: joint g177 (B4) @(-42, 1134) /w:[ 12 -1 11 18 ]
  //: joint g228 (B6) @(-1255, 1947) /w:[ 4 -1 3 26 ]
  assign B6 = B[6]; //: TAP g209 @(854,402) /sn:0 /R:2 /w:[ 15 3 4 ] /ss:0
  FA g96 (.b(w301), .a(w257), .Cin(w274), .Cout(w275), .S(w276));   //: @(-1608, 2117) /sz:(84, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g221 (A7) @(-1289, 1389) /w:[ -1 6 5 24 ]
  assign B5 = B[5]; //: TAP g196 @(854,383) /sn:0 /R:2 /w:[ 15 5 6 ] /ss:0
  NandAND g117 (.in2(A4), .in1(B7), .out(w5));   //: @(-1303, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>25 Bo0<0 ]
  FA g19 (.b(w62), .a(w21), .Cin(w50), .Cout(w52), .S(w55));   //: @(172, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g114 (.b(w5), .a(w294), .Cin(w329), .Cout(w330), .S(P11));   //: @(-1386, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g125 (B0) @(624, 295) /w:[ 12 -1 11 18 ]
  NandAND g78 (.in2(B4), .in1(A6), .out(w225));   //: @(-1090, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>25 Bo0<1 ]
  //: joint g223 (A0) @(-255, 1666) /w:[ -1 2 1 28 ]
  //: joint g219 (A5) @(-857, 1394) /w:[ -1 6 5 24 ]
  //: joint g155 (A7) @(-508, 88) /w:[ 14 -1 13 16 ]
  NandAND g113 (.in2(A7), .in1(B7), .out(w304));   //: @(-1928, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  FA g63 (.b(w199), .a(w202), .Cin(w176), .Cout(w161), .S(w177));   //: @(-368, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g93 (.b(w25), .a(w19), .Cin(w228), .Cout(w260), .S(w265));   //: @(-561, 1848) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g100 (.b(w286), .a(w252), .Cin(w287), .Cout(w288), .S(w289));   //: @(-1179, 2117) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g105 (.b(w280), .a(w247), .Cin(w302), .Cout(w287), .S(w303));   //: @(-997, 2117) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g244 (A2) @(-643, 1942) /w:[ -1 2 1 28 ]
  //: joint g215 (B5) @(-1041, 1674) /w:[ 4 -1 3 26 ]
  //: joint g212 (B5) @(-398, 1413) /w:[ 10 -1 9 20 ]
  //: joint g211 (A1) @(-263, 1399) /w:[ -1 4 3 26 ]
  //: joint g205 (A4) @(-443, 884) /w:[ -1 8 7 22 ]
  NandAND g101 (.in2(A0), .in1(B7), .out(w132));   //: @(-461, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>17 Bo0<1 ]
  FA g38 (.b(w70), .a(w22), .Cin(w60), .Cout(w114), .S(w31));   //: @(-14, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: IN g0 (A) @(857,245) /sn:0 /R:1 /w:[ 0 ]
  FA g43 (.b(w87), .a(w31), .Cin(w115), .Cout(w116), .S(w183));   //: @(-11, 1033) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  NandAND g48 (.in2(A3), .in1(B3), .out(w85));   //: @(-266, 892) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>23 Ti1>23 Bo0<0 ]
  //: joint g237 (B7) @(-614, 2211) /w:[ 12 -1 11 18 ]
  FA g37 (.b(w65), .a(w17), .Cin(w114), .Cout(w90), .S(w128));   //: @(-192, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  NandAND g122 (.in2(B7), .in1(A2), .out(w346));   //: @(-918, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  NandAND g120 (.in2(B7), .in1(A6), .out(w306));   //: @(-1694, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  NandAND g80 (.in2(B5), .in1(A1), .out(w224));   //: @(-277, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>27 Bo0<1 ]
  HA g95 (.b(w132), .a(w265), .Cout(w270), .S(P7));   //: @(-560, 2117) /sz:(72, 72) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<1 Bo0<0 ]
  FA g76 (.b(w217), .a(w172), .Cin(w191), .Cout(w214), .S(w4));   //: @(-1388, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g189 (B3) @(-627, 1130) /w:[ -1 4 3 26 ]
  //: joint g170 (A4) @(-269, 602) /w:[ -1 10 9 20 ]
  //: joint g152 (B2) @(-36, 612) /w:[ 8 -1 7 22 ]
  NandAND g75 (.in2(B4), .in1(A4), .out(w269));   //: @(-658, 1430) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>25 Bo0<1 ]
  assign A3 = A[3]; //: TAP g178 @(855,171) /sn:0 /R:2 /w:[ 15 7 8 ] /ss:0
  HA g44 (.b(w105), .a(w180), .Cout(w115), .S(P3));   //: @(187, 1033) /sz:(72, 72) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  assign B4 = B[4]; //: TAP g182 @(854,366) /sn:0 /R:2 /w:[ 15 7 8 ] /ss:0
  NandAND g16 (.in2(A6), .in1(B1), .out(w48));   //: @(-602, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>29 Bo0<0 ]
  NandAND g3 (.in2(A0), .in1(B0), .out(P0));   //: @(657, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>17 Bo0<0 ]
  assign A6 = A[6]; //: TAP g159 @(855,111) /sn:0 /R:2 /w:[ 15 13 14 ] /ss:0
  FA g47 (.b(w142), .a(w86), .Cin(w123), .Cout(w111), .S(w169));   //: @(-767, 1031) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g143 (B2) @(310, 612) /w:[ 12 -1 11 18 ]
  NandAND g26 (.in2(A2), .in1(B2), .out(w70));   //: @(98, 628) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>21 Bo0<0 ]
  FA g90 (.b(w8), .a(w214), .Cin(w233), .Cout(w256), .S(w257));   //: @(-1606, 1848) /sz:(87, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  HA g109 (.b(w350), .a(w307), .Cout(w312), .S(P8));   //: @(-754, 2371) /sz:(72, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  assign A1 = A[1]; //: TAP g158 @(855,204) /sn:0 /R:2 /w:[ 15 3 4 ] /ss:0
  HA g2 (.b(w49), .a(w0), .Cout(w2), .S(P1));   //: @(538, 512) /sz:(72, 72) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  //: joint g174 (A7) @(-662, 581) /w:[ -1 12 11 18 ]
  //: joint g128 (B0) @(450, 295) /w:[ 10 -1 9 20 ]
  FA g23 (.b(w24), .a(w45), .Cin(w59), .Cout(w6), .S(w37));   //: @(-374, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  FA g91 (.b(w20), .a(w205), .Cin(w260), .Cout(w245), .S(w261));   //: @(-765, 1848) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g141 (A6) @(-315, 111) /w:[ 14 -1 13 16 ]
  //: joint g127 (A1) @(594, 204) /w:[ 14 -1 13 16 ]
  NandAND g39 (.in2(A2), .in1(B3), .out(w92));   //: @(-82, 892) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>23 Ti1>21 Bo0<0 ]
  FA g24 (.b(w39), .a(w48), .Cin(w6), .Cout(w77), .S(w35));   //: @(-571, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g86 (.b(w18), .a(w63), .Cin(w245), .Cout(w246), .S(w247));   //: @(-996, 1848) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g104 (.b(w67), .a(w256), .Cin(w275), .Cout(w298), .S(w299));   //: @(-1805, 2117) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign P = {P15, P14, P13, P12, P11, P10, P9, P8, P7, P6, P5, P4, P3, P2, P1, P0}; //: CONCAT g250  @(851,2449) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  NandAND g29 (.in2(A7), .in1(B1), .out(w82));   //: @(-682, 629) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  FA g60 (.b(w211), .a(w169), .Cin(w162), .Cout(w148), .S(w241));   //: @(-766, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g110 (.b(w306), .a(w299), .Cin(w316), .Cout(w317), .S(P13));   //: @(-1812, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  FA g121 (.b(w346), .a(w303), .Cin(w312), .Cout(w344), .S(P9));   //: @(-992, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g168 (A2) @(118, 603) /w:[ -1 10 9 20 ]
  //: joint g248 (A6) @(-1468, 1935) /w:[ -1 2 1 28 ]
  //: joint g199 (A2) @(-245, 1121) /w:[ -1 6 5 24 ]
  NandAND g18 (.in2(A7), .in1(B0), .out(w39));   //: @(-528, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  FA g82 (.b(w11), .a(w4), .Cin(w232), .Cout(w233), .S(w234));   //: @(-1389, 1848) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g245 (A3) @(-846, 1942) /w:[ -1 2 1 28 ]
  NandAND g94 (.in2(B6), .in1(A1), .out(w25));   //: @(-451, 1690) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>29 Bo0<1 ]
  FA g119 (.b(w337), .a(w289), .Cin(w344), .Cout(w329), .S(P10));   //: @(-1181, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g173 (B2) @(-617, 876) /w:[ -1 2 1 28 ]
  //: joint g166 (A0) @(482, 603) /w:[ -1 10 9 20 ]
  //: joint g154 (A5) @(-385, 132) /w:[ 12 -1 11 18 ]
  FA g107 (.b(w140), .a(w261), .Cin(w270), .Cout(w302), .S(w307));   //: @(-764, 2117) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g216 (B5) @(-1265, 1674) /w:[ 2 -1 1 28 ]
  //: joint g188 (B3) @(-413, 876) /w:[ 6 -1 5 24 ]
  //: joint g184 (A0) @(302, 870) /w:[ -1 8 7 22 ]
  //: joint g172 (B2) @(-409, 612) /w:[ 4 -1 3 26 ]
  //: joint g193 (A7) @(-828, 839) /w:[ -1 10 9 20 ]
  FA g50 (.b(w85), .a(w93), .Cin(w136), .Cout(w122), .S(w202));   //: @(-368, 1031) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g133 (B1) @(189, 312) /w:[ 10 -1 9 20 ]
  NandAND g73 (.in2(A0), .in1(B5), .out(w262));   //: @(-89, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>17 Bo0<1 ]
  NandAND g9 (.in2(A4), .in1(B0), .out(w30));   //: @(26, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>25 Bo0<0 ]
  FA g68 (.b(w225), .a(w220), .Cin(w190), .Cout(w191), .S(w16));   //: @(-1185, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g225 (B6) @(-613, 1947) /w:[ -1 10 9 20 ]
  //: joint g186 (A2) @(-62, 870) /w:[ -1 8 7 22 ]
  //: joint g169 (A3) @(-66, 605) /w:[ -1 10 9 20 ]
  NandAND g71 (.in2(A7), .in1(B4), .out(w217));   //: @(-1309, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<1 ]
  NandAND g59 (.in2(A0), .in1(B4), .out(w189));   //: @(100, 1149) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>17 Bo0<0 ]
  FA g31 (.b(w58), .a(w55), .Cin(w56), .Cout(w60), .S(w180));   //: @(178, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  FA g22 (.b(w33), .a(w36), .Cin(w9), .Cout(w59), .S(w17));   //: @(-199, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g102 (.b(w291), .a(w234), .Cin(w288), .Cout(w274), .S(w294));   //: @(-1389, 2117) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g249 (A7) @(-1671, 1931) /w:[ -1 2 1 28 ]
  //: joint g231 (A3) @(-638, 1682) /w:[ -1 4 3 26 ]
  NandAND g87 (.in2(B6), .in1(A0), .out(w28));   //: @(-269, 1692) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>29 Bo0<1 ]
  //: joint g180 (B4) @(150, 1134) /w:[ 14 -1 13 16 ]
  NandAND g99 (.in2(A7), .in1(B6), .out(w67));   //: @(-1691, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  NandAND g83 (.in2(B5), .in1(A3), .out(w20));   //: @(-652, 1693) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>23 Ti1>27 Bo0<1 ]
  //: joint g203 (B4) @(-1046, 1411) /w:[ 2 -1 1 28 ]
  NandAND g41 (.in2(A7), .in1(B2), .out(w144));   //: @(-848, 892) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<1 ]
  FA g36 (.b(w73), .a(w37), .Cin(w90), .Cout(w74), .S(w93));   //: @(-371, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA g45 (.b(w135), .a(w78), .Cin(w122), .Cout(w123), .S(w124));   //: @(-563, 1031) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g213 (B5) @(-608, 1674) /w:[ -1 8 7 22 ]
  //: joint g156 (B1) @(-552, 312) /w:[ 2 -1 1 28 ]
  //: joint g138 (B1) @(-178, 312) /w:[ 6 -1 5 24 ]
  NandAND g69 (.in2(A2), .in1(B5), .out(w264));   //: @(-448, 1429) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>21 Bo0<1 ]
  FA g42 (.b(w144), .a(w110), .Cin(w111), .Cout(w94), .S(w157));   //: @(-978, 1031) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g167 (A1) @(280, 602) /w:[ -1 10 9 20 ]
  //: joint g151 (A4) @(-208, 149) /w:[ 12 -1 11 18 ]
  NandAND g66 (.in2(B4), .in1(A1), .out(w185));   //: @(-86, 1144) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>25 Bo0<0 ]
  //: joint g233 (A5) @(-1071, 1667) /w:[ -1 4 3 26 ]
  //: joint g232 (A4) @(-850, 1667) /w:[ -1 4 3 26 ]
  //: joint g191 (A5) @(-439, 602) /w:[ -1 10 9 20 ]
  //: joint g162 (B3) @(-32, 876) /w:[ 10 -1 9 20 ]
  //: joint g153 (B2) @(-239, 612) /w:[ 6 -1 5 24 ]
  //: joint g146 (B2) @(512, 612) /w:[ 14 -1 13 16 ]
  //: joint g242 (B7) @(-1650, 2211) /w:[ 2 -1 1 28 ]
  //: joint g241 (B7) @(-1438, 2211) /w:[ 4 -1 3 26 ]
  //: joint g239 (B7) @(-1031, 2211) /w:[ 8 -1 7 22 ]
  FA g34 (.b(w76), .a(w35), .Cin(w74), .Cout(w75), .S(w78));   //: @(-566, 781) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  NandAND g28 (.in2(A3), .in1(B2), .out(w65));   //: @(-86, 628) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>21 Ti1>23 Bo0<0 ]
  NandAND g46 (.in2(A0), .in1(B3), .out(w105));   //: @(282, 892) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>23 Ti1>17 Bo0<0 ]
  NandAND g57 (.in2(A7), .in1(B3), .out(w159));   //: @(-1083, 1150) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<0 ]
  FA g118 (.b(w304), .a(w298), .Cin(w317), .Cout(P15), .S(P14));   //: @(-2005, 2371) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  NandAND g11 (.in2(A3), .in1(B0), .out(w62));   //: @(217, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>23 Bo0<0 ]
  NandAND g14 (.in2(A6), .in1(B0), .out(w24));   //: @(-335, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>17 Ti1>29 Bo0<0 ]
  NandAND g84 (.in2(B5), .in1(A5), .out(w14));   //: @(-1085, 1690) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>27 Bo0<1 ]
  //: joint g5 (B0) @(707, 295) /w:[ 14 -1 13 16 ]
  //: joint g150 (A3) @(-31, 171) /w:[ 12 -1 11 18 ]
  //: joint g201 (B4) @(-614, 1411) /w:[ -1 6 5 24 ]
  NandAND g112 (.in2(B7), .in1(A5), .out(w335));   //: @(-1482, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  //: joint g187 (A3) @(-246, 870) /w:[ -1 8 7 22 ]
  FA g21 (.b(w30), .a(w42), .Cin(w52), .Cout(w9), .S(w22));   //: @(-18, 512) /sz:(82, 75) /sn:0 /anc:1 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  NandAND g61 (.in2(A3), .in1(B4), .out(w207));   //: @(-452, 1161) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>23 Bo0<0 ]
  //: joint g123 (A0) @(677, 225) /w:[ 14 -1 13 16 ]
  FA g79 (.b(w224), .a(w177), .Cin(w186), .Cout(w218), .S(w223));   //: @(-367, 1577) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  NandAND g20 (.in2(A5), .in1(B1), .out(w45));   //: @(-405, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>27 Bo0<0 ]
  NandAND g32 (.in2(B2), .in1(A5), .out(w76));   //: @(-453, 629) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>21 Bo0<0 ]
  NandAND g115 (.in2(A1), .in1(B7), .out(w350));   //: @(-664, 2224) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>19 Bo0<0 ]
  //: joint g240 (B7) @(-1253, 2211) /w:[ 6 -1 5 24 ]
  //: joint g235 (A7) @(-1478, 1640) /w:[ -1 4 3 26 ]
  assign A7 = A[7]; //: TAP g176 @(855,88) /sn:0 /R:2 /w:[ 15 15 16 ] /ss:0
  assign A2 = A[2]; //: TAP g175 @(855,189) /sn:0 /R:2 /w:[ 15 5 6 ] /ss:0
  NandAND g97 (.in2(A3), .in1(B6), .out(w280));   //: @(-866, 1960) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>29 Ti1>23 Bo0<0 ]
  //: joint g134 (B0) @(76, 295) /w:[ 6 -1 5 24 ]
  //: joint g145 (A0) @(516, 225) /w:[ 12 -1 11 18 ]
  //: joint g236 (B7) @(-411, 1942) /w:[ 14 -1 13 16 ]
  NandAND g15 (.in2(A3), .in1(B1), .out(w42));   //: @(-51, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>23 Bo0<0 ]
  NandAND g89 (.in2(A4), .in1(B5), .out(w18));   //: @(-870, 1689) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>27 Ti1>25 Bo0<1 ]
  //: joint g129 (A2) @(420, 189) /w:[ 14 -1 13 16 ]
  //: joint g148 (A1) @(347, 204) /w:[ 12 -1 11 18 ]
  //: joint g247 (A5) @(-1285, 1937) /w:[ -1 2 1 28 ]
  //: joint g227 (B6) @(-1037, 1947) /w:[ 6 -1 5 24 ]
  //: joint g202 (B4) @(-827, 1411) /w:[ 4 -1 3 26 ]
  assign B3 = B[3]; //: TAP g165 @(854,350) /sn:0 /R:2 /w:[ 15 9 10 ] /ss:0
  NandAND g27 (.in2(B2), .in1(A1), .out(w58));   //: @(266, 624) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>21 Bo0<0 ]
  assign B2 = B[2]; //: TAP g147 @(854,331) /sn:0 /R:2 /w:[ 15 11 12 ] /ss:0
  //: joint g218 (A4) @(-644, 1403) /w:[ -1 6 5 24 ]
  //: joint g171 (A6) @(-582, 290) /w:[ -1 12 11 18 ]
  assign B0 = B[0]; //: TAP g160 @(854,295) /sn:0 /R:2 /w:[ 15 15 16 ] /ss:0
  FA g62 (.b(w159), .a(w94), .Cin(w149), .Cout(w172), .S(w220));   //: @(-1184, 1295) /sz:(82, 75) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g238 (B7) @(-874, 2211) /w:[ 10 -1 9 20 ]
  //: joint g195 (B5) @(-39, 1413) /w:[ 14 -1 13 16 ]
  FA g88 (.b(w14), .a(w16), .Cin(w246), .Cout(w232), .S(w252));   //: @(-1184, 1848) /sz:(82, 75) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  NandAND g55 (.in2(A2), .in1(B4), .out(w199));   //: @(-265, 1150) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>25 Ti1>21 Bo0<0 ]
  //: joint g207 (A5) @(-657, 1120) /w:[ -1 8 7 22 ]
  HA g53 (.b(w189), .a(w183), .Cout(w145), .S(P4));   //: @(-10, 1295) /sz:(80, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  NandAND g13 (.in2(A4), .in1(B1), .out(w36));   //: @(-228, 341) /sz:(64, 93) /R:3 /sn:0 /p:[ Ti0>19 Ti1>25 Bo0<0 ]
  //: joint g135 (A4) @(46, 149) /w:[ 14 -1 13 16 ]
  //: joint g139 (A5) @(-134, 132) /w:[ 14 -1 13 16 ]
  //: joint g140 (B0) @(-285, 295) /w:[ 2 -1 1 28 ]

endmodule
//: /netlistEnd

//: /netlistBegin NandNOT
module NandNOT(out, in1);
//: interface  /sz:(93, 48) /bd:[ Li0>in1(16/48) Ro0<out(16/48) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(201,162)(201,214){1}
//: {2}(201,218)(201,270){3}
//: {4}(199,216)(170,216)(170,270){5}
output out;    //: /sn:0 {0}(201,359)(201,414){1}
//: enddecls

  //: comment g4 @(90,43) /sn:0
  //: /line:"La porta NOT si traduce in logica NAND come:"
  //: /line:""
  //: /line:" a' = (aa)'"
  //: /end
  //: joint g3 (in1) @(201, 216) /w:[ 2 -1 1 4 ]
  //: OUT g2 (out) @(201,411) /sn:0 /R:3 /w:[ 1 ]
  //: IN g1 (in1) @(201,160) /sn:0 /R:3 /w:[ 0 ]
  MyNAND g0 (.in1(in1), .in2(in1), .out(out));   //: @(153, 271) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>3 Ti1>5 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FS
module FS(PrIn, B, A, PrOut, D);
//: interface  /sz:(113, 44) /bd:[ Ti0>B(74/113) Ti1>A(36/113) Ri0>PrIn(16/44) Lo0<PrOut(22/44) Bo0<D(53/113) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(338,-67)(338,-40)(338,-40)(338,-12){1}
input PrIn;    //: /sn:0 {0}(379,-67)(379,117)(358,117)(358,168){1}
input A;    //: /sn:0 {0}(303,-67)(303,-37)(303,-37)(303,-12){1}
output PrOut;    //: /sn:0 {0}(245,349)(245,370)(245,370)(245,388){1}
output D;    //: /sn:0 {0}(345,282)(345,333)(345,333)(345,388){1}
wire w6;    //: /sn:0 {0}(262,260)(262,226)(305,226){1}
wire w3;    //: /sn:0 {0}(324,102)(324,168){1}
wire w2;    //: /sn:0 {0}(284,46)(225,46)(225,260){1}
//: enddecls

  //: IN g4 (PrIn) @(379,-69) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (B) @(338,-69) /sn:0 /R:3 /w:[ 0 ]
  HS g2 (.A(w3), .B(PrIn), .Pr(w6), .D(D));   //: @(306, 169) /sz:(74, 112) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  //: IN g1 (A) @(303,-69) /sn:0 /R:3 /w:[ 0 ]
  NandOR g6 (.in1(w6), .in2(w2), .out(PrOut));   //: @(209, 261) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<0 ]
  //: OUT g7 (PrOut) @(245,385) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g5 (D) @(345,385) /sn:0 /R:3 /w:[ 1 ]
  HS g0 (.A(A), .B(B), .Pr(w2), .D(w3));   //: @(285, -11) /sz:(75, 112) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin POT2
module POT2(P, F);
//: interface  /sz:(83, 74) /bd:[ Ti0>F[7:0](37/83) Bo0<P[15:0](40/83) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] F;    //: /sn:0 {0}(#:485,153)(485,119)(461,119){1}
//: {2}(459,117)(#:459,89){3}
//: {4}(457,119)(421,119)(#:421,153){5}
output [15:0] P;    //: /sn:0 {0}(#:458,255)(458,283)(459,283)(459,312){1}
//: enddecls

  //: OUT g3 (P) @(459,309) /sn:0 /R:3 /w:[ 1 ]
  //: joint g2 (F) @(459, 119) /w:[ 1 2 4 -1 ]
  //: IN g1 (F) @(459,87) /sn:0 /R:3 /w:[ 3 ]
  MUL16 g0 (.A(F), .B(F), .P(P));   //: @(403, 154) /sz:(109, 100) /sn:0 /p:[ Ti0>5 Ti1>0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin NandAND
module NandAND(out, in2, in1);
//: interface  /sz:(93, 64) /bd:[ Li0>in2(44/64) Li1>in1(14/64) Ro0<out(27/64) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(151,243)(151,210)(192,210)(192,169){1}
output out;    //: /sn:0 {0}(134,511)(134,552){1}
input in2;    //: /sn:0 {0}(128,243)(128,207)(84,207)(84,167){1}
wire w0;    //: /sn:0 {0}(136,331)(136,392){1}
//: {2}(138,394)(151,394)(151,422){3}
//: {4}(134,394)(119,394)(119,422){5}
//: enddecls

  MyNAND g4 (.in1(w0), .in2(w0), .out(out));   //: @(104, 423) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>3 Ti1>5 Bo0<0 ]
  //: OUT g2 (out) @(134,549) /sn:0 /R:3 /w:[ 1 ]
  //: IN g1 (in2) @(84,165) /sn:0 /R:3 /w:[ 1 ]
  MyNAND g6 (.in1(in1), .in2(in2), .out(w0));   //: @(106, 244) /sz:(60, 86) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  //: joint g5 (w0) @(136, 394) /w:[ 2 1 4 -1 ]
  //: IN g0 (in1) @(192,167) /sn:0 /R:3 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin HA
module HA(Cout, b, a, S);
//: interface  /sz:(72, 72) /bd:[ Ti0>a(18/72) Ti1>b(54/72) Lo0<Cout(33/72) Bo0<S(36/72) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(135,266)(135,204)(224,204){1}
//: {2}(226,206)(226,264){3}
//: {4}(226,202)(226,175){5}
output Cout;    //: /sn:0 {0}(142,406)(142,367){1}
input a;    //: /sn:0 {0}(151,266)(151,224)(260,224){1}
//: {2}(262,226)(262,264){3}
//: {4}(262,222)(262,173){5}
output S;    //: /sn:0 {0}(243,412)(243,365){1}
//: enddecls

  //: comment g4 @(58,-55) /sn:0
  //: /line:"L' Half Adder (HA) non prevede il riporto in ingresso, ma solo in uscita"
  //: /line:""
  //: /line:"La sua tabella di verità è:"
  //: /line:""
  //: /line:"  a | b | S | Cin"
  //: /line:" -----------------"
  //: /line:"  0 | 0 | 0 | 0"
  //: /line:"  0 | 1 | 1 | 0"
  //: /line:"  1 | 0 | 1 | 0"
  //: /line:"  1 | 1 | 0 | 1"
  //: /end
  //: OUT g8 (Cout) @(142,403) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (b) @(226,173) /sn:0 /R:3 /w:[ 5 ]
  //: IN g2 (a) @(262,171) /sn:0 /R:3 /w:[ 5 ]
  //: OUT g1 (S) @(243,409) /sn:0 /R:3 /w:[ 0 ]
  //: joint g6 (a) @(262, 224) /w:[ 2 -1 4 1 ]
  //: joint g7 (b) @(226, 204) /w:[ 2 -1 4 1 ]
  NandAND g5 (.in2(b), .in1(a), .out(Cout));   //: @(104, 267) /sz:(63, 99) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  NandEXOR g0 (.in1(a), .in2(b), .out(S));   //: @(207, 265) /sz:(64, 99) /R:3 /sn:0 /p:[ Ti0>3 Ti1>3 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FD16
module FD16(B, R, A, Q);
//: interface  /sz:(70, 54) /bd:[ Li0>A[15:0](10/54) Li1>B[15:0](38/54) Bo0<R[15:0](35/70) Ro0<Q[15:0](26/54) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [15:0] A;    //: /sn:0 {0}(#:1272,-297)(1262,-297)(1262,-297)(1258,-297){1}
//: {2}(1257,-297)(1237,-297){3}
//: {4}(1236,-297)(1212,-297){5}
//: {6}(1211,-297)(1186,-297){7}
//: {8}(1185,-297)(1163,-297){9}
//: {10}(1162,-297)(1142,-297){11}
//: {12}(1141,-297)(1121,-297){13}
//: {14}(1120,-297)(1101,-297){15}
//: {16}(1100,-297)(1082,-297){17}
//: {18}(1081,-297)(1064,-297){19}
//: {20}(1063,-297)(1047,-297){21}
//: {22}(1046,-297)(1027,-297){23}
//: {24}(1026,-297)(1008,-297){25}
//: {26}(1007,-297)(990,-297){27}
//: {28}(989,-297)(972,-297){29}
//: {30}(971,-297)(955,-297){31}
//: {32}(#:954,-297)(903,-297){33}
input [15:0] B;    //: /sn:0 {0}(#:862,-298)(837,-298){1}
//: {2}(836,-298)(819,-298){3}
//: {4}(818,-298)(797,-298){5}
//: {6}(796,-298)(775,-298){7}
//: {8}(774,-298)(753,-298){9}
//: {10}(752,-298)(733,-298){11}
//: {12}(732,-298)(712,-298){13}
//: {14}(711,-298)(688,-298){15}
//: {16}(687,-298)(665,-298){17}
//: {18}(664,-298)(640,-298){19}
//: {20}(639,-298)(615,-298){21}
//: {22}(614,-298)(588,-298){23}
//: {24}(587,-298)(561,-298){25}
//: {26}(560,-298)(534,-298){27}
//: {28}(533,-298)(507,-298){29}
//: {30}(506,-298)(481,-298){31}
//: {32}(#:480,-298)(427,-298){33}
output [15:0] Q;    //: /sn:0 {0}(4167,2507)(4135,2507)(4135,2507)(#:4101,2507){1}
supply0 w1444;    //: /sn:0 {0}(-1751,157)(-1751,131){1}
//: {2}(-1749,129)(-1571,129){3}
//: {4}(-1567,129)(-1387,129){5}
//: {6}(-1383,129)(-1205,129){7}
//: {8}(-1201,129)(-1023,129){9}
//: {10}(-1019,129)(-839,129){11}
//: {12}(-835,129)(-655,129){13}
//: {14}(-651,129)(-470,129){15}
//: {16}(-466,129)(-285,129){17}
//: {18}(-281,129)(-101,129){19}
//: {20}(-97,129)(87,129){21}
//: {22}(91,129)(267,129){23}
//: {24}(271,129)(451,129){25}
//: {26}(455,129)(618,129){27}
//: {28}(622,129)(928,129)(928,188){29}
//: {30}(930,190)(1099,190)(1099,361){31}
//: {32}(1101,363)(1278,363)(1278,527){33}
//: {34}(1280,529)(1453,529)(1453,690){35}
//: {36}(1455,692)(1634,692)(1634,859){37}
//: {38}(1636,861)(1819,861)(1819,1029){39}
//: {40}(1821,1031)(2018,1031)(2018,1188){41}
//: {42}(2020,1190)(2204,1190)(2204,1346){43}
//: {44}(2206,1348)(2371,1348)(2371,1498){45}
//: {46}(2373,1500)(2564,1500)(2564,1645){47}
//: {48}(2566,1647)(2763,1647)(2763,1798){49}
//: {50}(2765,1800)(2955,1800)(2955,1949){51}
//: {52}(2957,1951)(3122,1951)(3122,2100){53}
//: {54}(3124,2102)(3310,2102)(3310,2248){55}
//: {56}(3312,2250)(3496,2250)(3496,2402){57}
//: {58}(3498,2404)(3667,2404)(3667,2548){59}
//: {60}(3669,2550)(3705,2550)(3705,2556){61}
//: {62}(3665,2550)(3650,2550){63}
//: {64}(3494,2404)(3463,2404){65}
//: {66}(3308,2250)(3270,2250){67}
//: {68}(3120,2102)(3086,2102){69}
//: {70}(2953,1951)(2902,1951){71}
//: {72}(2761,1800)(2713,1800){73}
//: {74}(2562,1647)(2518,1647){75}
//: {76}(2369,1500)(2332,1500){77}
//: {78}(2202,1348)(2155,1348){79}
//: {80}(2016,1190)(1979,1190){81}
//: {82}(1817,1031)(1785,1031){83}
//: {84}(1632,861)(1591,861){85}
//: {86}(1451,692)(1411,692){87}
//: {88}(1276,529)(1229,529){89}
//: {90}(1097,363)(1058,363){91}
//: {92}(926,190)(882,190){93}
//: {94}(620,131)(620,157){95}
//: {96}(453,131)(453,157){97}
//: {98}(269,131)(269,157){99}
//: {100}(89,131)(-25:89,157){101}
//: {102}(-99,131)(-99,157){103}
//: {104}(-283,131)(-283,157){105}
//: {106}(-468,131)(-468,157){107}
//: {108}(-653,131)(-25:-653,157){109}
//: {110}(-837,131)(-837,157){111}
//: {112}(-1021,131)(-1021,157){113}
//: {114}(-1203,131)(-1203,157){115}
//: {116}(-1385,131)(-25:-1385,157){117}
//: {118}(-1569,131)(-1569,157){119}
//: {120}(-1753,129)(-1935,129)(-1935,157){121}
output [15:0] R;    //: /sn:0 {0}(4167,2758)(4134,2758)(4134,2758)(#:4106,2758){1}
wire w1049;    //: /sn:0 {0}(327,1719)(327,1747)(494,1747)(24:494,1767){1}
wire w471;    //: /sn:0 {0}(1024,933)(1024,968)(1184,968)(62:1184,998){1}
wire w457;    //: /sn:0 {0}(-835,933)(-835,998){1}
wire w864;    //: /sn:0 {0}(1145,1614)(1145,1572){1}
wire w602;    //: /sn:0 {0}(43:1740,1315)(1740,1290)(1559,1290)(1559,1262){1}
wire w605;    //: /sn:0 {0}(-926,1240)(-926,1260)(-894,1260)(-894,1225)(-873,1225){1}
wire w1243;    //: /sn:0 {0}(24:1013,2217)(1013,2198)(854,2198)(854,2174){1}
wire w382;    //: /sn:0 {0}(271,601)(271,659){1}
wire w374;    //: /sn:0 {0}(798,601)(798,659){1}
wire w534;    //: /sn:0 {0}(271,933)(-25:271,998){1}
wire B5;    //: {0}(35:-58,157)(-58,-57)(733,-57)(733,-294){1}
wire w1474;    //: /sn:0 {0}(2155,2550)(2210,2550){1}
wire w1274;    //: /sn:0 {0}(2870,2322)(2870,2352)(3041,2352)(43:3041,2371){1}
wire w4;    //: /sn:0 {0}(-2049,176)(-2049,159)(-1999,159)(-1999,191)(-1971,191){1}
wire w1535;    //: /sn:0 {0}(2486,2622)(2486,2632){1}
wire w1310;    //: /sn:0 {0}(2248,2217)(2248,2174){1}
wire Cr29;    //: /sn:0 {0}(3463,2436)(3773,2436)(3773,2572)(4095,2572){1}
wire w1100;    //: /sn:0 {0}(2071,2069)(2071,2023){1}
wire w539;    //: /sn:0 {0}(-45,1103)(-45,1135)(130,1135)(43:130,1157){1}
wire w661;    //: /sn:0 {0}(1195,1103)(1195,1135)(1366,1135)(62:1366,1157){1}
wire w721;    //: /sn:0 {0}(-13,1349)(53,1349){1}
wire w1369;    //: /sn:0 {0}(2964,2404)(2902,2404){1}
wire w733;    //: /sn:0 {0}(30:1184,1315)(1184,1293)(1029,1293)(1029,1262){1}
wire w1512;    //: /sn:0 {0}(1200,2622)(1200,2632){1}
wire w1309;    //: /sn:0 {0}(30:2287,2217)(2287,2200)(2126,2200)(2126,2174){1}
wire w327;    //: /sn:0 {0}(622,601)(-25:622,659){1}
wire Cr17;    //: /sn:0 {0}(2155,1380)(3861,1380)(3861,2502)(4095,2502){1}
wire w716;    //: /sn:0 {0}(1327,1467)(1327,1420){1}
wire w1278;    //: /sn:0 {0}(62:1934,2217)(1934,2201)(1751,2201)(1751,2174){1}
wire w1235;    //: /sn:0 {0}(43:661,2217)(661,2198)(507,2198)(507,2174){1}
wire w196;    //: /sn:0 {0}(-1665,398)(-1605,398){1}
wire w42;    //: /sn:0 {0}(-596,435)(-596,474)(-427,474)(30:-427,496){1}
wire A2;    //: {0}(1:3182,2217)(3182,-220)(1212,-220)(1212,-293){1}
wire w1525;    //: /sn:0 {0}(62:3041,2517)(3041,2500)(2868,2500)(2868,2476){1}
wire w1385;    //: /sn:0 {0}(2713,2404)(2780,2404){1}
wire w190;    //: /sn:0 {0}(-1239,398)(-1299,398){1}
wire w680;    //: /sn:0 {0}(30:494,1315)(494,1292)(326,1292)(326,1262){1}
wire w775;    //: /sn:0 {0}(2248,1572)(2248,1614){1}
wire w905;    //: /sn:0 {0}(1785,1647)(1857,1647){1}
wire w1280;    //: /sn:0 {0}(1785,2282)(1857,2282){1}
wire w583;    //: /sn:0 {0}(1895,1262)(1895,1315){1}
wire w629;    //: /sn:0 {0}(327,1103)(327,1135)(494,1135)(24:494,1157){1}
wire w752;    //: /sn:0 {0}(-567,1383)(-504,1383){1}
wire w848;    //: /sn:0 {0}(-382,1535)(-319,1535){1}
wire w622;    //: /sn:0 {0}(-231,1103)(-231,1136)(-58,1136)(62:-58,1157){1}
wire w1315;    //: /sn:0 {0}(30:837,2217)(837,2199)(677,2199)(677,2174){1}
wire w559;    //: /sn:0 {0}(-1019,1103)(-1019,1118){1}
wire w690;    //: /sn:0 {0}(1785,1380)(1857,1380){1}
wire w1226;    //: /sn:0 {0}(760,2137)(706,2137){1}
wire w199;    //: /sn:0 {0}(-1515,435)(-1515,471)(-1344,471)(43:-1344,496){1}
wire w909;    //: /sn:0 {0}(1785,1679)(1857,1679){1}
wire w1420;    //: /sn:0 {0}(622,2322)(622,2371){1}
wire w1300;    //: /sn:0 {0}(1229,2285)(1289,2285){1}
wire w1126;    //: /sn:0 {0}(539,1954)(584,1954){1}
wire w1042;    //: /sn:0 {0}(91,1767)(91,1719){1}
wire Cr13;    //: /sn:0 {0}(1785,1063)(3887,1063)(3887,2482)(4095,2482){1}
wire w116;    //: /sn:0 {0}(-42,262)(-42,310)(130,310)(30:130,330){1}
wire w32;    //: /sn:0 {0}(-1019,330)(-1019,262){1}
wire w846;    //: /sn:0 {0}(62:-242,1614)(-242,1595)(-416,1595)(-416,1572){1}
wire w53;    //: /sn:0 {0}(-1862,349)(-1862,332)(-1815,332)(-1815,364)(-1787,364){1}
wire w528;    //: /sn:0 {0}(-135,1034)(-197,1034){1}
wire w1347;    //: /sn:0 {0}(3341,2436)(3270,2436){1}
wire w710;    //: /sn:0 {0}(24:1366,1315)(1366,1292)(1201,1292)(1201,1262){1}
wire w760;    //: /sn:0 {0}(-25:1507,1467)(1507,1420){1}
wire w89;    //: /sn:0 {0}(3270,2282)(3784,2282)(3784,2562)(4095,2562){1}
wire w469;    //: /sn:0 {0}(848,764)(848,807)(1013,807)(62:1013,828){1}
wire w445;    //: /sn:0 {0}(510,764)(510,806)(661,806)(30:661,828){1}
wire w392;    //: /sn:0 {0}(-226,764)(-226,803)(-58,803)(30:-58,828){1}
wire w615;    //: /sn:0 {0}(-25:1145,1157)(1145,1103){1}
wire w774;    //: /sn:0 {0}(2304,1572)(2304,1595)(2473,1595)(24:2473,1614){1}
wire w892;    //: /sn:0 {0}(-367,1634)(-367,1617)(-336,1617)(-336,1648)(-319,1648){1}
wire w336;    //: /sn:0 {0}(-504,695)(-567,695){1}
wire w263;    //: /sn:0 {0}(-1239,532)(-1299,532){1}
wire w167;    //: /sn:0 {0}(233,395)(175,395){1}
wire w664;    //: /sn:0 {0}(1327,1262)(-25:1327,1315){1}
wire w346;    //: /sn:0 {0}(-466,601)(-466,659){1}
wire w135;    //: /sn:0 {0}(62:-1710,330)(-1710,294)(-1883,294)(-1883,262){1}
wire w169;    //: /sn:0 {0}(327,435)(327,476)(494,476)(24:494,496){1}
wire w777;    //: /sn:0 {0}(622,1420)(622,1467){1}
wire w942;    //: /sn:0 {0}(-231,1719)(-231,1749)(-58,1749)(62:-58,1767){1}
wire w11;    //: /sn:0 {0}(584,190)(539,190){1}
wire w120;    //: /sn:0 {0}(-382,222)(-323,222)(-323,222)(-319,222){1}
wire w78;    //: /sn:0 {0}(882,561)(936,561){1}
wire w743;    //: /sn:0 {0}(-319,1351)(-382,1351){1}
wire B9;    //: {0}(24:-793,157)(-793,-164)(640,-164)(640,-294){1}
wire w1510;    //: /sn:0 {0}(1229,2553)(1289,2553){1}
wire w1482;    //: /sn:0 {0}(2713,2550)(2780,2550){1}
wire w339;    //: /sn:0 {0}(-25:-651,828)(-651,764){1}
wire w412;    //: /sn:0 {0}(-1317,850)(-1317,833)(-1284,833)(-1284,862)(-1239,862){1}
wire w1152;    //: /sn:0 {0}(1701,2069)(1701,2023){1}
wire w1053;    //: /sn:0 {0}(1379,1719)(1379,1749)(1546,1749)(43:1546,1767){1}
wire w500;    //: /sn:0 {0}(1562,1103)(1562,1136)(1740,1136)(30:1740,1157){1}
wire w896;    //: /sn:0 {0}(1058,1679)(1107,1679){1}
wire w43;    //: /sn:0 {0}(-651,496)(-651,435){1}
wire w1071;    //: /sn:0 {0}(1289,1983)(1229,1983){1}
wire w954;    //: /sn:0 {0}(-25:271,1614)(271,1572){1}
wire w1477;    //: /sn:0 {0}(2332,2582)(2396,2582){1}
wire w1426;    //: /sn:0 {0}(798,2322)(798,2371){1}
wire w538;    //: /sn:0 {0}(-97,933)(-97,998){1}
wire w603;    //: /sn:0 {0}(1507,1262)(1507,1315){1}
wire w961;    //: /sn:0 {0}(2490,1719)(2490,1752)(2668,1752)(24:2668,1767){1}
wire w1497;    //: /sn:0 {0}(43:1740,2517)(1740,2503)(1559,2503)(1559,2476){1}
wire w1231;    //: /sn:0 {0}(271,2174)(271,2189){1}
wire w344;    //: /sn:0 {0}(-97,764)(-97,828){1}
wire w1096;    //: /sn:0 {0}(2033,1983)(1979,1983){1}
wire w569;    //: /sn:0 {0}(24:-427,998)(-427,974)(-595,974)(-595,933){1}
wire w584;    //: /sn:0 {0}(146,1103)(146,1135)(310,1135)(30:310,1157){1}
wire w704;    //: /sn:0 {0}(706,1380)(760,1380){1}
wire w1390;    //: /sn:0 {0}(1195,2322)(1195,2353)(1366,2353)(62:1366,2371){1}
wire w1098;    //: /sn:0 {0}(1979,1951)(2033,1951){1}
wire w677;    //: /sn:0 {0}(1979,1348)(2033,1348){1}
wire w744;    //: /sn:0 {0}(-226,1420)(-226,1451)(-58,1451)(30:-58,1467){1}
wire w186;    //: /sn:0 {0}(-1299,366)(-1239,366){1}
wire w685;    //: /sn:0 {0}(510,1420)(510,1448)(661,1448)(30:661,1467){1}
wire w1204;    //: /sn:0 {0}(1058,2137)(1107,2137){1}
wire w1065;    //: /sn:0 {0}(1145,1918)(1145,1872){1}
wire w142;    //: /sn:0 {0}(-1327,262)(-1327,303)(-1162,303)(24:-1162,330){1}
wire w1507;    //: /sn:0 {0}(30:1184,2517)(1184,2502)(1029,2502)(1029,2476){1}
wire w1020;    //: /sn:0 {0}(798,1918)(798,1872){1}
wire w487;    //: /sn:0 {0}(1701,1157)(1701,1103){1}
wire w1488;    //: /sn:0 {0}(1663,2553)(1591,2553){1}
wire w1331;    //: /sn:0 {0}(674,2322)(674,2349)(837,2349)(43:837,2371){1}
wire w1212;    //: /sn:0 {0}(1145,2217)(1145,2174){1}
wire w1014;    //: /sn:0 {0}(-25:1145,1767)(1145,1719){1}
wire w470;    //: /sn:0 {0}(974,828)(974,764){1}
wire w148;    //: /sn:0 {0}(-1512,262)(-1512,302)(-1344,302)(30:-1344,330){1}
wire w370;    //: /sn:0 {0}(-1201,601)(-1201,659){1}
wire w156;    //: /sn:0 {0}(-1860,413)(-1860,433)(-1814,433)(-1814,398)(-1787,398){1}
wire w862;    //: /sn:0 {0}(1145,1420)(1145,1467){1}
wire w255;    //: /sn:0 {0}(175,561)(233,561){1}
wire w800;    //: /sn:0 {0}(882,1532)(936,1532){1}
wire w395;    //: /sn:0 {0}(-13,861)(53,861){1}
wire w308;    //: /sn:0 {0}(1327,764)(1327,828){1}
wire w573;    //: /sn:0 {0}(507,933)(507,971)(661,971)(43:661,998){1}
wire w654;    //: /sn:0 {0}(62:-612,1315)(-612,1293)(-785,1293)(-785,1262){1}
wire w856;    //: /sn:0 {0}(1701,1572)(-25:1701,1614){1}
wire w1486;    //: /sn:0 {0}(62:1546,2517)(1546,2503)(1377,2503)(1377,2476){1}
wire w1284;    //: /sn:0 {0}(-25:1895,2371)(1895,2322){1}
wire w1317;    //: /sn:0 {0}(706,2285)(760,2285){1}
wire w121;    //: /sn:0 {0}(-319,190)(-323,190)(-323,190)(-382,190){1}
wire w1466;    //: /sn:0 {0}(3238,2622)(3238,2632){1}
wire w1276;    //: /sn:0 {0}(368,2235)(368,2218)(399,2218)(399,2251)(417,2251){1}
wire w1150;    //: /sn:0 {0}(1701,1872)(1701,1918){1}
wire w1470;    //: /sn:0 {0}(62:2287,2517)(2287,2500)(2121,2500)(2121,2476){1}
wire w1370;    //: /sn:0 {0}(43:3225,2517)(3225,2499)(3054,2499)(3054,2476){1}
wire w1244;    //: /sn:0 {0}(798,2217)(798,2174){1}
wire w1191;    //: /sn:0 {0}(-25:2248,2069)(2248,2023){1}
wire w390;    //: /sn:0 {0}(1563,933)(1563,968)(1740,968)(24:1740,998){1}
wire w873;    //: /sn:0 {0}(798,1614)(798,1572){1}
wire w1237;    //: /sn:0 {0}(2298,2023)(2298,2054)(2473,2054)(62:2473,2069){1}
wire w1155;    //: /sn:0 {0}(2964,2134)(2902,2134){1}
wire Cr3;    //: /sn:0 {0}(882,222)(3981,222)(3981,2432)(4095,2432){1}
wire w935;    //: /sn:0 {0}(53,1650)(-13,1650){1}
wire w1338;    //: /sn:0 {0}(-25:974,2217)(974,2174){1}
wire w391;    //: /sn:0 {0}(1507,933)(1507,998){1}
wire w1319;    //: /sn:0 {0}(760,2253)(706,2253){1}
wire w1170;    //: /sn:0 {0}(2713,2134)(2780,2134){1}
wire w1412;    //: /sn:0 {0}(974,2322)(974,2371){1}
wire w1045;    //: /sn:0 {0}(1945,1719)(1945,1751)(2110,1751)(62:2110,1767){1}
wire w1029;    //: /sn:0 {0}(175,1835)(233,1835){1}
wire w1004;    //: /sn:0 {0}(1895,1918)(1895,1872){1}
wire w576;    //: /sn:0 {0}(622,1157)(622,1103){1}
wire w69;    //: /sn:0 {0}(1058,529)(1107,529){1}
wire w984;    //: /sn:0 {0}(2155,1832)(2210,1832){1}
wire w300;    //: /sn:0 {0}(-319,692)(-382,692){1}
wire w799;    //: /sn:0 {0}(974,1420)(974,1467){1}
wire w1508;    //: /sn:0 {0}(1145,2517)(1145,2476){1}
wire w1043;    //: /sn:0 {0}(43:310,1918)(310,1901)(143,1901)(143,1872){1}
wire w377;    //: /sn:0 {0}(-963,601)(-963,644)(-796,644)(24:-796,659){1}
wire w47;    //: /sn:0 {0}(853,435)(853,474)(1013,474)(30:1013,496){1}
wire w579;    //: /sn:0 {0}(1857,1222)(1785,1222){1}
wire w634;    //: /sn:0 {0}(91,1103)(91,1157){1}
wire w1421;    //: /sn:0 {0}(760,2407)(709,2407){1}
wire w1119;    //: /sn:0 {0}(1785,1983)(1857,1983){1}
wire w582;    //: /sn:0 {0}(1951,1262)(1951,1286)(2110,1286)(24:2110,1315){1}
wire w397;    //: /sn:0 {0}(30:130,998)(130,972)(-42,972)(-42,933){1}
wire w550;    //: /sn:0 {0}(-567,1034)(-504,1034){1}
wire w137;    //: /sn:0 {0}(-1849,225)(-1816,225)(-1816,225)(-1787,225){1}
wire w38;    //: /sn:0 {0}(974,496)(974,435){1}
wire w1122;    //: /sn:0 {0}(1895,2069)(1895,2023){1}
wire w107;    //: /sn:0 {0}(53,222)(-13,222){1}
wire w221;    //: /sn:0 {0}(-1676,579)(-1676,599)(-1632,599)(-1632,564)(-1605,564){1}
wire w1485;    //: /sn:0 {0}(2902,2582)(2964,2582){1}
wire w1105;    //: /sn:0 {0}(706,1952)(760,1952){1}
wire Cr9;    //: /sn:0 {0}(1411,724)(3918,724)(3918,2462)(4095,2462){1}
wire w724;    //: /sn:0 {0}(175,1383)(233,1383){1}
wire w1351;    //: /sn:0 {0}(3379,2476)(3379,2517){1}
wire w843;    //: /sn:0 {0}(-601,1420)(-601,1448)(-427,1448)(62:-427,1467){1}
wire w483;    //: /sn:0 {0}(1663,1063)(1591,1063){1}
wire w699;    //: /sn:0 {0}(1701,1467)(1701,1420){1}
wire w740;    //: /sn:0 {0}(-281,1262)(-281,1315){1}
wire w762;    //: /sn:0 {0}(-97,1262)(-25:-97,1315){1}
wire w1414;    //: /sn:0 {0}(1058,2407)(1107,2407){1}
wire w1238;    //: /sn:0 {0}(2434,2069)(2434,2023){1}
wire w491;    //: /sn:0 {0}(175,1031)(233,1031){1}
wire w745;    //: /sn:0 {0}(-281,1420)(-281,1467){1}
wire w891;    //: /sn:0 {0}(2071,1767)(2071,1719){1}
wire w1393;    //: /sn:0 {0}(1229,2405)(1289,2405){1}
wire w1372;    //: /sn:0 {0}(523,2391)(523,2380)(560,2380)(560,2405)(587,2405){1}
wire w1021;    //: /sn:0 {0}(1562,1719)(1562,1749)(1740,1749)(30:1740,1767){1}
wire w343;    //: /sn:0 {0}(-41,764)(-41,804)(130,804)(24:130,828){1}
wire w81;    //: /sn:0 {0}(974,601)(974,659){1}
wire w669;    //: /sn:0 {0}(674,1103)(674,1136)(837,1136)(43:837,1157){1}
wire w1517;    //: /sn:0 {0}(936,2553)(882,2553){1}
wire w1062;    //: /sn:0 {0}(2874,2023)(2874,2055)(3041,2055)(24:3041,2069){1}
wire w746;    //: /sn:0 {0}(-135,1383)(-197,1383){1}
wire B15;    //: {0}(18:-1894,157)(-1894,-269)(481,-269)(481,-294){1}
wire w1171;    //: /sn:0 {0}(2780,2102)(2713,2102){1}
wire w827;    //: /sn:0 {0}(43:661,1614)(661,1598)(507,1598)(507,1572){1}
wire w985;    //: /sn:0 {0}(2210,1800)(2155,1800){1}
wire w883;    //: /sn:0 {0}(2210,1647)(2155,1647){1}
wire w1059;    //: /sn:0 {0}(2780,1983)(2713,1983){1}
wire w22;    //: /sn:0 {0}(-935,222)(-873,222){1}
wire w495;    //: /sn:0 {0}(233,1063)(175,1063){1}
wire w1536;    //: /sn:0 {0}(4100,2743)(2434,2743)(2434,2622){1}
wire w1335;    //: /sn:0 {0}(2679,2322)(2679,2353)(2857,2353)(62:2857,2371){1}
wire w1106;    //: /sn:0 {0}(848,2023)(848,2051)(1013,2051)(62:1013,2069){1}
wire w122;    //: /sn:0 {0}(-229,262)(-229,310)(-58,310)(43:-58,330){1}
wire w1288;    //: /sn:0 {0}(2396,2282)(2332,2282){1}
wire w1511;    //: /sn:0 {0}(1107,2553)(1058,2553){1}
wire w1491;    //: /sn:0 {0}(4100,2793)(1507,2793)(1507,2622){1}
wire w1383;    //: /sn:0 {0}(-25:2629,2371)(2629,2322){1}
wire w1287;    //: /sn:0 {0}(-25:2434,2217)(2434,2174){1}
wire w917;    //: /sn:0 {0}(24:1013,1614)(1013,1599)(854,1599)(854,1572){1}
wire B2;    //: {0}(47:494,157)(494,15)(797,15)(797,-294){1}
wire w313;    //: /sn:0 {0}(936,692)(882,692){1}
wire w871;    //: /sn:0 {0}(2434,1767)(2434,1719){1}
wire w1120;    //: /sn:0 {0}(1857,1951)(1785,1951){1}
wire w442;    //: /sn:0 {0}(-281,828)(-281,764){1}
wire w335;    //: /sn:0 {0}(-651,601)(-651,659){1}
wire w701;    //: /sn:0 {0}(-747,1400)(-747,1420)(-716,1420)(-716,1383)(-689,1383){1}
wire w922;    //: /sn:0 {0}(622,1614)(622,1572){1}
wire w956;    //: /sn:0 {0}(271,1767)(271,1719){1}
wire Cr28;    //: /sn:0 {0}(882,2137)(936,2137){1}
wire w684;    //: /sn:0 {0}(417,1348)(355,1348){1}
wire w1263;    //: /sn:0 {0}(1663,2282)(1591,2282){1}
wire w1055;    //: /sn:0 {0}(43:1740,1918)(1740,1900)(1559,1900)(1559,1872){1}
wire w372;    //: /sn:0 {0}(-1201,764)(-1201,828){1}
wire w982;    //: /sn:0 {0}(2123,1719)(2123,1750)(2287,1750)(43:2287,1767){1}
wire Cr4;    //: /sn:0 {0}(1058,395)(3956,395)(3956,2442)(4095,2442){1}
wire w1375;    //: /sn:0 {0}(2071,2322)(2071,2371){1}
wire w801;    //: /sn:0 {0}(1107,1500)(1058,1500){1}
wire w1361;    //: /sn:0 {0}(3184,2371)(3184,2322){1}
wire w1182;    //: /sn:0 {0}(1557,2023)(1557,2049)(1740,2049)(62:1740,2069){1}
wire w1109;    //: /sn:0 {0}(24:1366,1918)(1366,1904)(1201,1904)(1201,1872){1}
wire w1031;    //: /sn:0 {0}(233,1803)(175,1803){1}
wire w503;    //: /sn:0 {0}(1327,933)(1327,998){1}
wire w545;    //: /sn:0 {0}(853,1103)(853,1136)(1013,1136)(30:1013,1157){1}
wire w586;    //: /sn:0 {0}(175,1222)(233,1222){1}
wire w803;    //: /sn:0 {0}(62:1184,1614)(1184,1597)(1024,1597)(1024,1572){1}
wire w841;    //: /sn:0 {0}(-97,1614)(-97,1572){1}
wire B8;    //: {0}(27:-612,157)(-612,-142)(665,-142)(665,-294){1}
wire w508;    //: /sn:0 {0}(-1126,1018)(-1126,1001)(-1085,1001)(-1085,1032)(-1057,1032){1}
wire w1289;    //: /sn:0 {0}(2518,2250)(2591,2250){1}
wire w1018;    //: /sn:0 {0}(798,1767)(798,1719){1}
wire w41;    //: /sn:0 {0}(-689,363)(-751,363){1}
wire w543;    //: /sn:0 {0}(706,1063)(760,1063){1}
wire w822;    //: /sn:0 {0}(-25:798,1467)(798,1420){1}
wire w1404;    //: /sn:0 {0}(1507,2517)(1507,2476){1}
wire Cr20;    //: /sn:0 {0}(175,1535)(233,1535){1}
wire w288;    //: /sn:0 {0}(91,601)(91,659){1}
wire w228;    //: /sn:0 {0}(-97,601)(-25:-97,659){1}
wire w847;    //: /sn:0 {0}(-466,1572)(-466,1587){1}
wire w926;    //: /sn:0 {0}(1507,1572)(1507,1614){1}
wire w1239;    //: /sn:0 {0}(62:2668,2217)(2668,2201)(2484,2201)(2484,2174){1}
wire B0;    //: {0}(15:837,157)(837,-294){1}
wire w1410;    //: /sn:0 {0}(2434,2517)(2434,2476){1}
wire w1132;    //: /sn:0 {0}(91,1918)(91,1872){1}
wire w1199;    //: /sn:0 {0}(974,2069)(974,2023){1}
wire w1037;    //: /sn:0 {0}(53,1803)(-13,1803){1}
wire w1032;    //: /sn:0 {0}(30:494,1918)(494,1900)(326,1900)(326,1872){1}
wire w279;    //: /sn:0 {0}(672,601)(672,638)(837,638)(62:837,659){1}
wire w1437;    //: /sn:0 {0}(2123,2322)(2123,2355)(2287,2355)(43:2287,2371){1}
wire w433;    //: /sn:0 {0}(-567,862)(-504,862){1}
wire w65;    //: /sn:0 {0}(505,435)(505,475)(661,475)(62:661,496){1}
wire A5;    //: {0}(2:2627,1767)(2627,-149)(1142,-149)(1142,-293){1}
wire w769;    //: /sn:0 {0}(2127,1420)(2127,1452)(2287,1452)(24:2287,1467){1}
wire w1286;    //: /sn:0 {0}(24:2473,2217)(2473,2200)(2304,2200)(2304,2174){1}
wire w1093;    //: /sn:0 {0}(1591,1983)(1663,1983){1}
wire w253;    //: /sn:0 {0}(146,435)(146,472)(310,472)(30:310,496){1}
wire w655;    //: /sn:0 {0}(-835,1262)(-835,1277){1}
wire w1134;    //: /sn:0 {0}(141,2023)(141,2049)(310,2049)(62:310,2069){1}
wire w348;    //: /sn:0 {0}(-466,828)(-466,764){1}
wire w825;    //: /sn:0 {0}(323,1420)(323,1449)(494,1449)(43:494,1467){1}
wire w1342;    //: /sn:0 {0}(2071,2217)(2071,2174){1}
wire w378;    //: /sn:0 {0}(-835,601)(-25:-835,659){1}
wire w1165;    //: /sn:0 {0}(30:1546,2217)(1546,2202)(1382,2202)(1382,2174){1}
wire w1115;    //: /sn:0 {0}(1026,2023)(1026,2050)(1184,2050)(43:1184,2069){1}
wire w480;    //: /sn:0 {0}(455,933)(455,998){1}
wire w784;    //: /sn:0 {0}(1950,1420)(1950,1451)(2110,1451)(30:2110,1467){1}
wire w831;    //: /sn:0 {0}(1229,1532)(1289,1532){1}
wire w1034;    //: /sn:0 {0}(417,1835)(355,1835){1}
wire w1033;    //: /sn:0 {0}(271,1918)(271,1872){1}
wire w225;    //: /sn:0 {0}(53,529)(-13,529){1}
wire w683;    //: /sn:0 {0}(539,1348)(584,1348){1}
wire w788;    //: /sn:0 {0}(30:2287,1614)(2287,1594)(2126,1594)(2126,1572){1}
wire w413;    //: /sn:0 {0}(-1315,914)(-1315,934)(-1283,934)(-1283,896)(-1239,896){1}
wire w234;    //: /sn:0 {0}(355,529)(417,529){1}
wire w1469;    //: /sn:0 {0}(685,2595)(685,2615)(726,2615)(726,2585)(757,2585){1}
wire w402;    //: /sn:0 {0}(1229,893)(1289,893){1}
wire w1128;    //: /sn:0 {0}(510,2023)(510,2051)(661,2051)(30:661,2069){1}
wire w766;    //: /sn:0 {0}(974,1262)(974,1315){1}
wire w270;    //: /sn:0 {0}(-1517,601)(-1517,645)(-1344,645)(62:-1344,659){1}
wire w23;    //: /sn:0 {0}(760,222)(706,222){1}
wire w70;    //: /sn:0 {0}(1201,601)(1201,636)(1366,636)(24:1366,659){1}
wire w84;    //: /sn:0 {0}(850,601)(850,638)(1013,638)(43:1013,659){1}
wire B11;    //: {0}(21:-1162,157)(-1162,-206)(588,-206)(588,-294){1}
wire w1057;    //: /sn:0 {0}(2685,1872)(2685,1900)(2857,1900)(24:2857,1918){1}
wire w24;    //: /sn:0 {0}(798,330)(798,262){1}
wire w566;    //: /sn:0 {0}(1145,933)(1145,998){1}
wire w1479;    //: /sn:0 {0}(-25:2818,2517)(2818,2476){1}
wire w1056;    //: /sn:0 {0}(1507,1872)(1507,1918){1}
wire w649;    //: /sn:0 {0}(-466,1262)(-466,1315){1}
wire w317;    //: /sn:0 {0}(-1486,742)(-1486,762)(-1448,762)(-1448,727)(-1421,727){1}
wire w1445;    //: /sn:0 {0}(3463,2550)(3528,2550){1}
wire w986;    //: /sn:0 {0}(43:2473,1918)(2473,1899)(2300,1899)(2300,1872){1}
wire w328;    //: /sn:0 {0}(584,724)(539,724){1}
wire w354;    //: /sn:0 {0}(455,828)(455,764){1}
wire w333;    //: /sn:0 {0}(706,724)(760,724){1}
wire w853;    //: /sn:0 {0}(1557,1420)(1557,1451)(1740,1451)(62:1740,1467){1}
wire w1396;    //: /sn:0 {0}(1411,2439)(1469,2439){1}
wire w330;    //: /sn:0 {0}(539,692)(584,692){1}
wire w925;    //: /sn:0 {0}(30:1546,1614)(1546,1596)(1382,1596)(1382,1572){1}
wire w1072;    //: /sn:0 {0}(30:2668,1918)(2668,1899)(2489,1899)(2489,1872){1}
wire w631;    //: /sn:0 {0}(24:661,1315)(661,1292)(511,1292)(511,1262){1}
wire w1428;    //: /sn:0 {0}(798,2476)(798,2517){1}
wire w422;    //: /sn:0 {0}(678,764)(678,806)(837,806)(24:837,828){1}
wire w670;    //: /sn:0 {0}(798,1157)(798,1103){1}
wire w773;    //: /sn:0 {0}(2155,1500)(2210,1500){1}
wire w920;    //: /sn:0 {0}(974,1767)(974,1719){1}
wire w461;    //: /sn:0 {0}(-1057,864)(-1117,864){1}
wire w432;    //: /sn:0 {0}(-319,864)(-382,864){1}
wire w332;    //: /sn:0 {0}(622,828)(622,764){1}
wire w763;    //: /sn:0 {0}(-41,1420)(-41,1452)(130,1452)(24:130,1467){1}
wire w394;    //: /sn:0 {0}(-197,893)(-135,893){1}
wire w1101;    //: /sn:0 {0}(2155,1983)(2210,1983){1}
wire w997;    //: /sn:0 {0}(1411,1832)(1469,1832){1}
wire w526;    //: /sn:0 {0}(62:-242,998)(-242,975)(-416,975)(-416,933){1}
wire w61;    //: /sn:0 {0}(-410,435)(-410,472)(-242,472)(24:-242,496){1}
wire w913;    //: /sn:0 {0}(355,1648)(417,1648){1}
wire w1380;    //: /sn:0 {0}(-25:2071,2517)(2071,2476){1}
wire w885;    //: /sn:0 {0}(2248,1767)(2248,1719){1}
wire w614;    //: /sn:0 {0}(1030,1103)(1030,1135)(1184,1135)(24:1184,1157){1}
wire w617;    //: /sn:0 {0}(1229,1190)(1289,1190){1}
wire Cr34;    //: /sn:0 {0}(1411,2585)(1469,2585){1}
wire w57;    //: /sn:0 {0}(-1117,364)(-1057,364){1}
wire w77;    //: /sn:0 {0}(-319,561)(-382,561){1}
wire A15;    //: {0}(796,157)(59:796,112)(955,112)(955,-293){1}
wire w778;    //: /sn:0 {0}(539,1532)(584,1532){1}
wire Cr10;    //: /sn:0 {0}(-751,727)(-689,727){1}
wire w58;    //: /sn:0 {0}(-969,435)(-969,473)(-796,473)(62:-796,496){1}
wire w240;    //: /sn:0 {0}(-689,532)(-751,532){1}
wire w1202;    //: /sn:0 {0}(62:1184,2217)(1184,2199)(1024,2199)(1024,2174){1}
wire w859;    //: /sn:0 {0}(24:310,1614)(310,1599)(147,1599)(147,1572){1}
wire w992;    //: /sn:0 {0}(1229,1832)(1289,1832){1}
wire w1054;    //: /sn:0 {0}(1507,1767)(1507,1719){1}
wire w1254;    //: /sn:0 {0}(24:3418,2371)(3418,2350)(3241,2350)(3241,2322){1}
wire w972;    //: /sn:0 {0}(936,1800)(882,1800){1}
wire w1117;    //: /sn:0 {0}(30:1934,1918)(1934,1902)(1756,1902)(1756,1872){1}
wire w620;    //: /sn:0 {0}(1145,1262)(1145,1315){1}
wire w987;    //: /sn:0 {0}(2248,1918)(2248,1872){1}
wire w1261;    //: /sn:0 {0}(1562,2322)(1562,2354)(1740,2354)(30:1740,2371){1}
wire w20;    //: /sn:0 {0}(1979,1222)(3876,1222)(3876,2492)(4095,2492){1}
wire w1181;    //: /sn:0 {0}(184,2153)(184,2173)(211,2173)(211,2137)(233,2137){1}
wire w261;    //: /sn:0 {0}(-1299,564)(-1239,564){1}
wire w515;    //: /sn:0 {0}(505,1103)(505,1135)(661,1135)(62:661,1157){1}
wire w1236;    //: /sn:0 {0}(455,2217)(455,2174){1}
wire w218;    //: /sn:0 {0}(798,496)(798,435){1}
wire w574;    //: /sn:0 {0}(622,933)(622,998){1}
wire w1334;    //: /sn:0 {0}(2629,2217)(2629,2174){1}
wire w639;    //: /sn:0 {0}(882,1222)(936,1222){1}
wire w952;    //: /sn:0 {0}(-25:1895,1767)(1895,1719){1}
wire w1019;    //: /sn:0 {0}(43:1013,1918)(1013,1902)(850,1902)(850,1872){1}
wire w409;    //: /sn:0 {0}(1107,861)(1058,861){1}
wire w1323;    //: /sn:0 {0}(62:494,2217)(494,2200)(321,2200)(321,2174){1}
wire w364;    //: /sn:0 {0}(-1383,601)(-1383,659){1}
wire w531;    //: /sn:0 {0}(-25:-281,1157)(-281,1103){1}
wire w360;    //: /sn:0 {0}(-964,764)(-964,805)(-796,805)(30:-796,828){1}
wire w247;    //: /sn:0 {0}(-225,601)(-225,642)(-58,642)(24:-58,659){1}
wire w590;    //: /sn:0 {0}(271,1262)(271,1315){1}
wire w594;    //: /sn:0 {0}(1591,1222)(1663,1222){1}
wire w665;    //: /sn:0 {0}(-410,1103)(-410,1136)(-242,1136)(24:-242,1157){1}
wire w719;    //: /sn:0 {0}(91,1262)(91,1315){1}
wire w555;    //: /sn:0 {0}(-1151,933)(-1151,975)(-980,975)(62:-980,998){1}
wire w635;    //: /sn:0 {0}(43:310,1315)(310,1291)(143,1291)(143,1262){1}
wire w911;    //: /sn:0 {0}(455,1614)(455,1572){1}
wire w1297;    //: /sn:0 {0}(1058,2251)(1107,2251){1}
wire w1163;    //: /sn:0 {0}(1411,2102)(1469,2102){1}
wire w459;    //: /sn:0 {0}(-1333,764)(-1333,803)(-1162,803)(62:-1162,828){1}
wire w919;    //: /sn:0 {0}(1030,1719)(1030,1749)(1184,1749)(24:1184,1767){1}
wire w426;    //: /sn:0 {0}(706,861)(760,861){1}
wire w630;    //: /sn:0 {0}(-25:455,1157)(455,1103){1}
wire w1136;    //: /sn:0 {0}(175,1986)(233,1986){1}
wire w115;    //: /sn:0 {0}(-135,190)(-133,190)(-133,190)(-197,190){1}
wire w1307;    //: /sn:0 {0}(1379,2322)(1379,2354)(1546,2354)(43:1546,2371){1}
wire w1484;    //: /sn:0 {0}(4100,2723)(2818,2723)(2818,2622){1}
wire w910;    //: /sn:0 {0}(62:494,1614)(494,1599)(321,1599)(321,1572){1}
wire w28;    //: /sn:0 {0}(854,262)(854,298)(1013,298)(24:1013,330){1}
wire w563;    //: /sn:0 {0}(-783,1103)(-783,1131)(-612,1131)(43:-612,1157){1}
wire w889;    //: /sn:0 {0}(2033,1647)(1979,1647){1}
wire w974;    //: /sn:0 {0}(974,1918)(974,1872){1}
wire w443;    //: /sn:0 {0}(43:-58,998)(-58,974)(-229,974)(-229,933){1}
wire w1175;    //: /sn:0 {0}(2629,2069)(2629,2023){1}
wire w1002;    //: /sn:0 {0}(1785,1800)(1857,1800){1}
wire w652;    //: /sn:0 {0}(-835,1103)(-835,1157){1}
wire w1185;    //: /sn:0 {0}(1857,2102)(1785,2102){1}
wire w1225;    //: /sn:0 {0}(622,2217)(622,2174){1}
wire w272;    //: /sn:0 {0}(-1483,564)(-1421,564){1}
wire w1521;    //: /sn:0 {0}(43:1013,2517)(1013,2500)(850,2500)(850,2476){1}
wire w1135;    //: /sn:0 {0}(91,2023)(91,2038){1}
wire w454;    //: /sn:0 {0}(-751,864)(-689,864){1}
wire w1480;    //: /sn:0 {0}(2780,2582)(2713,2582){1}
wire w1129;    //: /sn:0 {0}(455,2069)(455,2023){1}
wire w700;    //: /sn:0 {0}(-749,1336)(-749,1319)(-716,1319)(-716,1349)(-689,1349){1}
wire w805;    //: /sn:0 {0}(1058,1532)(1107,1532){1}
wire w1262;    //: /sn:0 {0}(1507,2371)(1507,2322){1}
wire w1365;    //: /sn:0 {0}(3186,2517)(3186,2476){1}
wire w6;    //: /sn:0 {0}(-1057,193)(-1063,193)(-1063,193)(-1117,193){1}
wire w522;    //: /sn:0 {0}(882,1031)(936,1031){1}
wire w485;    //: /sn:0 {0}(1591,1031)(1663,1031){1}
wire w7;    //: /sn:0 {0}(355,222)(417,222){1}
wire w314;    //: /sn:0 {0}(1026,764)(1026,805)(1184,805)(43:1184,828){1}
wire w34;    //: /sn:0 {0}(882,363)(936,363){1}
wire w552;    //: /sn:0 {0}(-596,1103)(-596,1133)(-427,1133)(30:-427,1157){1}
wire w1392;    //: /sn:0 {0}(1469,2407)(1411,2407){1}
wire w379;    //: /sn:0 {0}(-779,764)(-779,804)(-612,804)(24:-612,828){1}
wire w162;    //: /sn:0 {0}(-231,435)(-231,471)(-58,471)(62:-58,496){1}
wire w648;    //: /sn:0 {0}(30:-242,1315)(-242,1293)(-411,1293)(-411,1262){1}
wire w702;    //: /sn:0 {0}(62:837,1315)(837,1293)(672,1293)(672,1262){1}
wire w713;    //: /sn:0 {0}(1411,1348)(1469,1348){1}
wire w1320;    //: /sn:0 {0}(853,2322)(853,2351)(1013,2351)(30:1013,2371){1}
wire Cr24;    //: /sn:0 {0}(539,1835)(585,1835){1}
wire w322;    //: /sn:0 {0}(-13,692)(53,692){1}
wire w756;    //: /sn:0 {0}(-466,1420)(-466,1467){1}
wire w1409;    //: /sn:0 {0}(30:2668,2517)(2668,2502)(2489,2502)(2489,2476){1}
wire w1407;    //: /sn:0 {0}(2332,2436)(2396,2436){1}
wire w1312;    //: /sn:0 {0}(2210,2250)(2155,2250){1}
wire w1242;    //: /sn:0 {0}(-25:798,2069)(798,2023){1}
wire w1161;    //: /sn:0 {0}(1327,2023)(1327,2069){1}
wire w1158;    //: /sn:0 {0}(3058,2174)(3058,2200)(3224,2200)(24:3224,2217){1}
wire w427;    //: /sn:0 {0}(854,933)(854,968)(1013,968)(24:1013,998){1}
wire w1210;    //: /sn:0 {0}(1145,2069)(1145,2023){1}
wire w154;    //: /sn:0 {0}(-1749,262)(-1749,330){1}
wire w71;    //: /sn:0 {0}(1145,601)(1145,659){1}
wire Cr32;    //: /sn:0 {0}(1229,2439)(1289,2439){1}
wire w1292;    //: /sn:0 {0}(2434,2371)(2434,2322){1}
wire w1075;    //: /sn:0 {0}(2591,1951)(2518,1951){1}
wire w527;    //: /sn:0 {0}(-281,933)(-281,998){1}
wire w352;    //: /sn:0 {0}(417,692)(355,692){1}
wire w168;    //: /sn:0 {0}(175,363)(233,363){1}
wire w63;    //: /sn:0 {0}(-783,435)(-783,473)(-612,473)(43:-612,496){1}
wire w577;    //: /sn:0 {0}(1757,1103)(1757,1136)(1934,1136)(24:1934,1157){1}
wire w1074;    //: /sn:0 {0}(2518,1983)(2591,1983){1}
wire w623;    //: /sn:0 {0}(-97,1157)(-97,1103){1}
wire w650;    //: /sn:0 {0}(-319,1225)(-382,1225){1}
wire w789;    //: /sn:0 {0}(2071,1572)(2071,1614){1}
wire w1389;    //: /sn:0 {0}(2713,2436)(2780,2436){1}
wire w1006;    //: /sn:0 {0}(505,1719)(505,1748)(660,1748)(62:660,1767){1}
wire w1419;    //: /sn:0 {0}(505,2322)(505,2347)(664,2347)(62:664,2371){1}
wire w1374;    //: /sn:0 {0}(1945,2322)(1945,2354)(2110,2354)(62:2110,2371){1}
wire w596;    //: /sn:0 {0}(1756,1262)(1756,1288)(1934,1288)(30:1934,1315){1}
wire w829;    //: /sn:0 {0}(1200,1420)(1200,1450)(1366,1450)(30:1366,1467){1}
wire Cr21;    //: /sn:0 {0}(2518,1679)(3835,1679)(3835,2522)(4095,2522){1}
wire w1513;    //: /sn:0 {0}(4100,2813)(1145,2813)(1145,2622){1}
wire w1362;    //: /sn:0 {0}(3086,2436)(3148,2436){1}
wire w468;    //: /sn:0 {0}(-1019,933)(-1019,998){1}
wire w1458;    //: /sn:0 {0}(3270,2582)(3341,2582){1}
wire w463;    //: /sn:0 {0}(-1201,933)(-1201,948){1}
wire w224;    //: /sn:0 {0}(-197,561)(-135,561){1}
wire w863;    //: /sn:0 {0}(43:1366,1614)(1366,1597)(1197,1597)(1197,1572){1}
wire w916;    //: /sn:0 {0}(539,1682)(584,1682){1}
wire B10;    //: {0}(22:-980,157)(-980,-189)(615,-189)(615,-294){1}
wire w1504;    //: /sn:0 {0}(2591,2550)(2518,2550){1}
wire w741;    //: /sn:0 {0}(-382,1383)(-319,1383){1}
wire w244;    //: /sn:0 {0}(-751,564)(-689,564){1}
wire w193;    //: /sn:0 {0}(-1605,366)(-1665,366){1}
wire w581;    //: /sn:0 {0}(1785,1190)(1857,1190){1}
wire w1194;    //: /sn:0 {0}(2155,2102)(2210,2102){1}
wire w1173;    //: /sn:0 {0}(2818,2174)(2818,2217){1}
wire w597;    //: /sn:0 {0}(1701,1262)(1701,1315){1}
wire w681;    //: /sn:0 {0}(455,1262)(455,1315){1}
wire w696;    //: /sn:0 {0}(1591,1380)(1663,1380){1}
wire w1318;    //: /sn:0 {0}(882,2253)(936,2253){1}
wire w852;    //: /sn:0 {0}(-281,1572)(-281,1614){1}
wire w588;    //: /sn:0 {0}(233,1190)(175,1190){1}
wire w618;    //: /sn:0 {0}(1058,1190)(1107,1190){1}
wire w1011;    //: /sn:0 {0}(-25:622,1918)(622,1873){1}
wire w667;    //: /sn:0 {0}(24:-58,1315)(-58,1293)(-225,1293)(-225,1262){1}
wire w686;    //: /sn:0 {0}(455,1420)(455,1467){1}
wire A14;    //: {0}(11:972,330)(972,-293){1}
wire w419;    //: /sn:0 {0}(62:494,998)(494,970)(321,970)(321,933){1}
wire w505;    //: /sn:0 {0}(1289,1031)(1229,1031){1}
wire w811;    //: /sn:0 {0}(24:1740,1614)(1740,1597)(1564,1597)(1564,1572){1}
wire w1027;    //: /sn:0 {0}(146,1719)(146,1748)(310,1748)(30:310,1767){1}
wire w448;    //: /sn:0 {0}(584,861)(539,861){1}
wire w242;    //: /sn:0 {0}(-785,601)(-785,643)(-612,643)(62:-612,659){1}
wire w50;    //: /sn:0 {0}(584,363)(539,363){1}
wire w712;    //: /sn:0 {0}(1289,1380)(1229,1380){1}
wire w861;    //: /sn:0 {0}(1026,1420)(1026,1450)(1184,1450)(43:1184,1467){1}
wire w1509;    //: /sn:0 {0}(1058,2585)(1107,2585){1}
wire w39;    //: /sn:0 {0}(-751,395)(-689,395){1}
wire Cr14;    //: /sn:0 {0}(-382,1066)(-319,1066){1}
wire w663;    //: /sn:0 {0}(62:1546,1315)(1546,1292)(1377,1292)(1377,1262){1}
wire w783;    //: /sn:0 {0}(760,1532)(706,1532){1}
wire w876;    //: /sn:0 {0}(760,1647)(706,1647){1}
wire w323;    //: /sn:0 {0}(141,764)(141,805)(310,805)(62:310,828){1}
wire w3;    //: /sn:0 {0}(417,190)(355,190){1}
wire w1267;    //: /sn:0 {0}(2964,2250)(2902,2250){1}
wire Cr27;    //: /sn:0 {0}(3086,2134)(3798,2134)(3798,2552)(4095,2552){1}
wire w845;    //: /sn:0 {0}(-319,1503)(-382,1503){1}
wire w1391;    //: /sn:0 {0}(1327,2371)(1327,2322){1}
wire w29;    //: /sn:0 {0}(-595,262)(-595,308)(-427,308)(24:-427,330){1}
wire w30;    //: /sn:0 {0}(-780,262)(-780,309)(-612,309)(30:-612,330){1}
wire w817;    //: /sn:0 {0}(175,1501)(233,1501){1}
wire w351;    //: /sn:0 {0}(355,724)(417,724){1}
wire w651;    //: /sn:0 {0}(-969,1103)(-969,1131)(-796,1131)(62:-796,1157){1}
wire w915;    //: /sn:0 {0}(-25:455,1767)(455,1719){1}
wire w329;    //: /sn:0 {0}(706,692)(760,692){1}
wire w736;    //: /sn:0 {0}(1107,1348)(1058,1348){1}
wire B7;    //: {0}(29:-427,157)(-427,-113)(688,-113)(688,-294){1}
wire w1397;    //: /sn:0 {0}(1757,2322)(1757,2353)(1934,2353)(24:1934,2371){1}
wire w1272;    //: /sn:0 {0}(2713,2282)(2780,2282){1}
wire w851;    //: /sn:0 {0}(43:-58,1614)(-58,1597)(-229,1597)(-229,1572){1}
wire w507;    //: /sn:0 {0}(1327,1157)(1327,1103){1}
wire w489;    //: /sn:0 {0}(91,933)(91,998){1}
wire w1378;    //: /sn:0 {0}(1979,2404)(2033,2404){1}
wire w31;    //: /sn:0 {0}(-835,330)(-835,262){1}
wire w795;    //: /sn:0 {0}(1895,1572)(1895,1614){1}
wire w628;    //: /sn:0 {0}(-13,1225)(53,1225){1}
wire w266;    //: /sn:0 {0}(-1057,564)(-1117,564){1}
wire w821;    //: /sn:0 {0}(678,1420)(678,1449)(837,1449)(24:837,1467){1}
wire w1524;    //: /sn:0 {0}(4100,2823)(974,2823)(974,2622){1}
wire w1266;    //: /sn:0 {0}(2902,2282)(2964,2282){1}
wire w517;    //: /sn:0 {0}(539,1063)(584,1063){1}
wire w557;    //: /sn:0 {0}(-873,1034)(-935,1034){1}
wire A11;    //: {0}(7:1505,828)(1505,-13)(1027,-13)(1027,-293){1}
wire w521;    //: /sn:0 {0}(1058,1031)(1107,1031){1}
wire w428;    //: /sn:0 {0}(798,933)(798,998){1}
wire w1041;    //: /sn:0 {0}(-45,1719)(-45,1749)(130,1749)(43:130,1767){1}
wire w707;    //: /sn:0 {0}(848,1420)(848,1451)(1013,1451)(62:1013,1467){1}
wire w1430;    //: /sn:0 {0}(2818,2371)(2818,2322){1}
wire w67;    //: /sn:0 {0}(1107,561)(1058,561){1}
wire w1180;    //: /sn:0 {0}(183,2089)(183,2072)(213,2072)(213,2103)(233,2103){1}
wire w284;    //: /sn:0 {0}(-1019,601)(-1019,659){1}
wire w1456;    //: /sn:0 {0}(30:3418,2517)(3418,2496)(3241,2496)(3241,2476){1}
wire w1424;    //: /sn:0 {0}(709,2439)(760,2439){1}
wire w1520;    //: /sn:0 {0}(882,2585)(936,2585){1}
wire w1172;    //: /sn:0 {0}(2873,2174)(2873,2201)(3041,2201)(30:3041,2217){1}
wire B4;    //: {0}(37:130,157)(130,-36)(753,-36)(753,-294){1}
wire w1387;    //: /sn:0 {0}(24:2857,2517)(2857,2501)(2685,2501)(2685,2476){1}
wire w320;    //: /sn:0 {0}(-13,724)(53,724){1}
wire w726;    //: /sn:0 {0}(622,1262)(-25:622,1315){1}
wire w933;    //: /sn:0 {0}(-13,1682)(53,1682){1}
wire w1514;    //: /sn:0 {0}(1289,2585)(1229,2585){1}
wire w447;    //: /sn:0 {0}(539,893)(584,893){1}
wire w417;    //: /sn:0 {0}(417,861)(355,861){1}
wire w717;    //: /sn:0 {0}(1411,1380)(1469,1380){1}
wire w1221;    //: /sn:0 {0}(539,2137)(584,2137){1}
wire w399;    //: /sn:0 {0}(53,893)(-13,893){1}
wire w496;    //: /sn:0 {0}(1382,933)(1382,969)(1546,969)(30:1546,998){1}
wire w720;    //: /sn:0 {0}(233,1351)(175,1351){1}
wire w1443;    //: /sn:0 {0}(3528,2582)(3463,2582){1}
wire w291;    //: /sn:0 {0}(1289,724)(1229,724){1}
wire w1464;    //: /sn:0 {0}(3086,2582)(3148,2582){1}
wire w1377;    //: /sn:0 {0}(2210,2404)(2155,2404){1}
wire w358;    //: /sn:0 {0}(-935,695)(-873,695){1}
wire w72;    //: /sn:0 {0}(-567,561)(-504,561){1}
wire w948;    //: /sn:0 {0}(-97,1767)(-97,1719){1}
wire w1174;    //: /sn:0 {0}(2486,2023)(2486,2054)(2668,2054)(43:2668,2069){1}
wire w337;    //: /sn:0 {0}(-751,693)(-689,693){1}
wire w1423;    //: /sn:0 {0}(625,2476)(625,2491){1}
wire w1355;    //: /sn:0 {0}(1785,2404)(1857,2404){1}
wire w1251;    //: /sn:0 {0}(3146,2282)(3086,2282){1}
wire w117;    //: /sn:0 {0}(-97,330)(-97,262){1}
wire w159;    //: /sn:0 {0}(-382,395)(-319,395){1}
wire w1279;    //: /sn:0 {0}(1895,2217)(1895,2174){1}
wire w1257;    //: /sn:0 {0}(1507,2217)(1507,2174){1}
wire w1447;    //: /sn:0 {0}(4100,2683)(3566,2683)(3566,2622){1}
wire w1178;    //: /sn:0 {0}(43:2857,2217)(2857,2201)(2681,2201)(2681,2174){1}
wire w1040;    //: /sn:0 {0}(-13,1835)(53,1835){1}
wire w141;    //: /sn:0 {0}(-1483,193)(-1443,193)(-1443,193)(-1421,193){1}
wire w227;    //: /sn:0 {0}(-47,601)(-47,641)(130,641)(62:130,659){1}
wire w368;    //: /sn:0 {0}(-1299,727)(-1239,727){1}
wire w217;    //: /sn:0 {0}(674,435)(674,475)(837,475)(43:837,496){1}
wire w1527;    //: /sn:0 {0}(3052,2622)(3052,2631){1}
wire w1141;    //: /sn:0 {0}(62:2287,1918)(2287,1902)(2121,1902)(2121,1872){1}
wire w638;    //: /sn:0 {0}(974,1157)(974,1103){1}
wire A12;    //: {0}(7:1325,659)(1325,16)(1008,16)(1008,-293){1}
wire w1367;    //: /sn:0 {0}(3002,2371)(3002,2322){1}
wire w1245;    //: /sn:0 {0}(1753,2023)(1753,2050)(1934,2050)(43:1934,2069){1}
wire w355;    //: /sn:0 {0}(-1146,601)(-1146,643)(-980,643)(30:-980,659){1}
wire w1496;    //: /sn:0 {0}(4100,2763)(2071,2763)(2071,2622){1}
wire w456;    //: /sn:0 {0}(30:-612,998)(-612,975)(-780,975)(-780,933){1}
wire Cr7;    //: /sn:0 {0}(-1117,398)(-1057,398){1}
wire w816;    //: /sn:0 {0}(417,1503)(355,1503){1}
wire w449;    //: /sn:0 {0}(677,933)(677,970)(837,970)(30:837,998){1}
wire w1147;    //: /sn:0 {0}(678,2023)(678,2052)(837,2052)(24:837,2069){1}
wire w794;    //: /sn:0 {0}(43:2110,1614)(2110,1594)(1947,1594)(1947,1572){1}
wire w802;    //: /sn:0 {0}(882,1500)(936,1500){1}
wire w809;    //: /sn:0 {0}(1593,1500)(1663,1500){1}
wire w1438;    //: /sn:0 {0}(2248,2322)(2248,2371){1}
wire w1229;    //: /sn:0 {0}(417,2105)(355,2105){1}
wire w899;    //: /sn:0 {0}(1195,1719)(1195,1750)(1366,1750)(62:1366,1767){1}
wire w1515;    //: /sn:0 {0}(675,2476)(675,2502)(835,2502)(62:835,2517){1}
wire w840;    //: /sn:0 {0}(30:130,1614)(130,1597)(-42,1597)(-42,1572){1}
wire w779;    //: /sn:0 {0}(706,1500)(760,1500){1}
wire w1273;    //: /sn:0 {0}(2780,2250)(2713,2250){1}
wire w163;    //: /sn:0 {0}(-25:-281,496)(-281,435){1}
wire w1468;    //: /sn:0 {0}(683,2531)(683,2514)(728,2514)(728,2551)(757,2551){1}
wire w149;    //: /sn:0 {0}(-1567,262)(-1567,330){1}
wire w975;    //: /sn:0 {0}(1107,1832)(1058,1832){1}
wire w1166;    //: /sn:0 {0}(1327,2217)(1327,2174){1}
wire w326;    //: /sn:0 {0}(511,601)(511,638)(661,638)(24:661,659){1}
wire w5;    //: /sn:0 {0}(-25:272,330)(272,262){1}
wire w613;    //: /sn:0 {0}(706,1222)(760,1222){1}
wire w718;    //: /sn:0 {0}(-47,1262)(-47,1293)(130,1293)(62:130,1315){1}
wire w748;    //: /sn:0 {0}(-651,1262)(-651,1315){1}
wire w928;    //: /sn:0 {0}(1469,1647)(1411,1647){1}
wire w1069;    //: /sn:0 {0}(1200,2023)(1200,2049)(1366,2049)(30:1366,2069){1}
wire w600;    //: /sn:0 {0}(1411,1222)(1469,1222){1}
wire w1434;    //: /sn:0 {0}(1145,2322)(-25:1145,2371){1}
wire w1039;    //: /sn:0 {0}(-97,1872)(-97,1887){1}
wire Cr6;    //: /sn:0 {0}(-1299,225)(-1253,225)(-1253,225)(-1239,225){1}
wire w424;    //: /sn:0 {0}(760,893)(706,893){1}
wire w806;    //: /sn:0 {0}(1383,1420)(1383,1451)(1547,1451)(24:1547,1467){1}
wire w499;    //: /sn:0 {0}(1469,1031)(1411,1031){1}
wire w525;    //: /sn:0 {0}(1058,1063)(1107,1063){1}
wire w786;    //: /sn:0 {0}(1979,1532)(2033,1532){1}
wire w790;    //: /sn:0 {0}(1753,1420)(1753,1451)(1934,1451)(43:1934,1467){1}
wire w1505;    //: /sn:0 {0}(2684,2622)(2684,2632){1}
wire w438;    //: /sn:0 {0}(-25:91,828)(91,764){1}
wire w0;    //: /sn:0 {0}(1591,893)(3898,893)(3898,2472)(4095,2472){1}
wire w189;    //: /sn:0 {0}(-1383,496)(-1383,435){1}
wire w226;    //: /sn:0 {0}(-197,529)(-135,529){1}
wire w1094;    //: /sn:0 {0}(24:2110,1918)(2110,1902)(1951,1902)(1951,1872){1}
wire w549;    //: /sn:0 {0}(-751,1066)(-689,1066){1}
wire A6;    //: {0}(2:2432,1614)(2432,-126)(1121,-126)(1121,-293){1}
wire w1190;    //: /sn:0 {0}(2127,2023)(2127,2053)(2287,2053)(24:2287,2069){1}
wire w403;    //: /sn:0 {0}(1289,861)(1229,861){1}
wire w1523;    //: /sn:0 {0}(1026,2622)(1026,2632){1}
wire w1313;    //: /sn:0 {0}(30:2473,2371)(2473,2356)(2303,2356)(2303,2322){1}
wire w1073;    //: /sn:0 {0}(2629,1872)(2629,1918){1}
wire w19;    //: /sn:0 {0}(706,190)(760,190){1}
wire w12;    //: /sn:0 {0}(-873,190)(-935,190){1}
wire w501;    //: /sn:0 {0}(1507,1157)(1507,1103){1}
wire w714;    //: /sn:0 {0}(1229,1348)(1289,1348){1}
wire w1167;    //: /sn:0 {0}(1469,2134)(1411,2134){1}
wire w570;    //: /sn:0 {0}(-466,933)(-25:-466,998){1}
wire w1304;    //: /sn:0 {0}(1701,2371)(1701,2322){1}
wire w1528;    //: /sn:0 {0}(4100,2713)(3002,2713)(3002,2622){1}
wire w104;    //: /sn:0 {0}(-2047,240)(-2047,260)(-1998,260)(-1998,225)(-1971,225){1}
wire w838;    //: /sn:0 {0}(-13,1503)(53,1503){1}
wire w872;    //: /sn:0 {0}(30:837,1614)(837,1598)(677,1598)(677,1572){1}
wire w551;    //: /sn:0 {0}(-689,1034)(-751,1034){1}
wire w1492;    //: /sn:0 {0}(1591,2585)(1663,2585){1}
wire w1460;    //: /sn:0 {0}(3434,2622)(3434,2632){1}
wire B6;    //: {0}(31:-242,157)(-242,-88)(712,-88)(712,-294){1}
wire w1454;    //: /sn:0 {0}(4100,2773)(1895,2773)(1895,2622){1}
wire w1408;    //: /sn:0 {0}(2396,2404)(2332,2404){1}
wire w1211;    //: /sn:0 {0}(43:1366,2217)(1366,2201)(1197,2201)(1197,2174){1}
wire w924;    //: /sn:0 {0}(622,1767)(622,1719){1}
wire w1451;    //: /sn:0 {0}(1979,2550)(2033,2550){1}
wire w1415;    //: /sn:0 {0}(936,2407)(882,2407){1}
wire w338;    //: /sn:0 {0}(-601,764)(-601,803)(-427,803)(62:-427,828){1}
wire w187;    //: /sn:0 {0}(-1421,366)(-1483,366){1}
wire w1373;    //: /sn:0 {0}(525,2455)(525,2467)(557,2467)(557,2439)(587,2439){1}
wire w1189;    //: /sn:0 {0}(1785,2134)(1857,2134){1}
wire w296;    //: /sn:0 {0}(-411,601)(-411,641)(-242,641)(30:-242,659){1}
wire w2;    //: /sn:0 {0}(175,222)(233,222){1}
wire w814;    //: /sn:0 {0}(141,1420)(141,1451)(310,1451)(62:310,1467){1}
wire w1399;    //: /sn:0 {0}(24:2110,2517)(2110,2499)(1951,2499)(1951,2476){1}
wire w1228;    //: /sn:0 {0}(271,2069)(271,2023){1}
wire w502;    //: /sn:0 {0}(1197,933)(1197,968)(1366,968)(43:1366,998){1}
wire w1449;    //: /sn:0 {0}(1895,2517)(1895,2476){1}
wire w554;    //: /sn:0 {0}(-504,1066)(-567,1066){1}
wire w785;    //: /sn:0 {0}(2071,1467)(2071,1420){1}
wire w1207;    //: /sn:0 {0}(24:1740,2217)(1740,2203)(1563,2203)(1563,2174){1}
wire w286;    //: /sn:0 {0}(91,435)(91,496){1}
wire w1386;    //: /sn:0 {0}(2518,2404)(2591,2404){1}
wire w1005;    //: /sn:0 {0}(1979,1832)(2033,1832){1}
wire w345;    //: /sn:0 {0}(-599,601)(-599,642)(-427,642)(43:-427,659){1}
wire w40;    //: /sn:0 {0}(-567,363)(-504,363){1}
wire w262;    //: /sn:0 {0}(-1117,532)(-1057,532){1}
wire w723;    //: /sn:0 {0}(91,1420)(-25:91,1467){1}
wire w1010;    //: /sn:0 {0}(62:837,1918)(837,1899)(672,1899)(672,1873){1}
wire w834;    //: /sn:0 {0}(1327,1614)(1327,1572){1}
wire w898;    //: /sn:0 {0}(1058,1647)(1107,1647){1}
wire w1518;    //: /sn:0 {0}(847,2622)(847,2631){1}
wire w1290;    //: /sn:0 {0}(2332,2250)(2396,2250){1}
wire w429;    //: /sn:0 {0}(882,893)(936,893){1}
wire w879;    //: /sn:0 {0}(936,1679)(882,1679){1}
wire w205;    //: /sn:0 {0}(-1145,435)(-1145,472)(-980,472)(24:-980,496){1}
wire w995;    //: /sn:0 {0}(62:1546,1918)(1546,1901)(1377,1901)(1377,1872){1}
wire w62;    //: /sn:0 {0}(-466,496)(-466,435){1}
wire w1322;    //: /sn:0 {0}(936,2285)(882,2285){1}
wire w241;    //: /sn:0 {0}(-935,530)(-873,530){1}
wire w897;    //: /sn:0 {0}(1289,1647)(1229,1647){1}
wire w82;    //: /sn:0 {0}(706,561)(760,561){1}
wire w519;    //: /sn:0 {0}(974,933)(-25:974,998){1}
wire Cr23;    //: /sn:0 {0}(2902,1983)(3814,1983)(3814,2542)(4095,2542){1}
wire w1339;    //: /sn:0 {0}(1030,2322)(1030,2352)(1184,2352)(24:1184,2371){1}
wire w452;    //: /sn:0 {0}(-835,764)(-835,828){1}
wire w37;    //: /sn:0 {0}(1030,435)(1030,470)(1184,470)(24:1184,496){1}
wire w170;    //: /sn:0 {0}(271,435)(271,496){1}
wire w625;    //: /sn:0 {0}(-197,1191)(-135,1191){1}
wire w751;    //: /sn:0 {0}(-651,1420)(-651,1435){1}
wire w1253;    //: /sn:0 {0}(3086,2250)(3146,2250){1}
wire w1223;    //: /sn:0 {0}(584,2105)(539,2105){1}
wire w1030;    //: /sn:0 {0}(355,1803)(417,1803){1}
wire w732;    //: /sn:0 {0}(271,1420)(271,1467){1}
wire w1133;    //: /sn:0 {0}(233,1954)(175,1954){1}
wire w21;    //: /sn:0 {0}(-751,190)(-689,190){1}
wire A9;    //: {0}(3:1893,1157)(1893,-59)(1064,-59)(1064,-293){1}
wire w561;    //: /sn:0 {0}(43:-796,998)(-796,974)(-967,974)(-967,933){1}
wire w927;    //: /sn:0 {0}(1411,1679)(1469,1679){1}
wire w293;    //: /sn:0 {0}(1229,692)(1289,692){1}
wire w1017;    //: /sn:0 {0}(674,1719)(674,1746)(837,1746)(43:837,1767){1}
wire w304;    //: /sn:0 {0}(1029,601)(1029,637)(1184,637)(30:1184,659){1}
wire w595;    //: /sn:0 {0}(1663,1190)(1591,1190){1}
wire w943;    //: /sn:0 {0}(-281,1719)(-281,1734){1}
wire w1476;    //: /sn:0 {0}(4100,2753)(2248,2753)(2248,2622){1}
wire w1104;    //: /sn:0 {0}(936,1954)(882,1954){1}
wire w316;    //: /sn:0 {0}(-1488,678)(-1488,661)(-1449,661)(-1449,693)(-1421,693){1}
wire w52;    //: /sn:0 {0}(622,496)(622,435){1}
wire w232;    //: /sn:0 {0}(417,561)(355,561){1}
wire w808;    //: /sn:0 {0}(1469,1532)(1411,1532){1}
wire w932;    //: /sn:0 {0}(91,1572)(91,1614){1}
wire w1452;    //: /sn:0 {0}(1857,2550)(1785,2550){1}
wire w1354;    //: /sn:0 {0}(1591,2436)(1663,2436){1}
wire w1184;    //: /sn:0 {0}(1591,2134)(1663,2134){1}
wire Cr12;    //: /sn:0 {0}(-567,896)(-504,896){1}
wire w991;    //: /sn:0 {0}(1327,1767)(1327,1719){1}
wire w400;    //: /sn:0 {0}(1200,764)(1200,806)(1366,806)(30:1366,828){1}
wire w146;    //: /sn:0 {0}(-1665,225)(-1629,225)(-1629,225)(-1605,225){1}
wire w1356;    //: /sn:0 {0}(1663,2404)(1591,2404){1}
wire w294;    //: /sn:0 {0}(1383,764)(1383,807)(1546,807)(24:1546,828){1}
wire w1296;    //: /sn:0 {0}(1289,2253)(1229,2253){1}
wire w297;    //: /sn:0 {0}(-281,601)(-281,659){1}
wire w161;    //: /sn:0 {0}(-382,363)(-319,363){1}
wire w506;    //: /sn:0 {0}(1379,1103)(1379,1136)(1546,1136)(43:1546,1157){1}
wire B3;    //: {0}(41:310,157)(310,-9)(775,-9)(775,-294){1}
wire w1530;    //: /sn:0 {0}(-25:1327,2517)(1327,2476){1}
wire w1473;    //: /sn:0 {0}(2396,2550)(2332,2550){1}
wire w653;    //: /sn:0 {0}(-689,1193)(-751,1193){1}
wire w703;    //: /sn:0 {0}(798,1262)(798,1315){1}
wire A4;    //: {0}(2:2816,1918)(2816,-175)(1163,-175)(1163,-293){1}
wire w1111;    //: /sn:0 {0}(1383,2023)(1383,2049)(1546,2049)(24:1546,2069){1}
wire w9;    //: /sn:0 {0}(175,190)(233,190){1}
wire w780;    //: /sn:0 {0}(584,1500)(539,1500){1}
wire w1095;    //: /sn:0 {0}(-25:2071,1918)(2071,1872){1}
wire w16;    //: /sn:0 {0}(455,330)(455,262){1}
wire w1282;    //: /sn:0 {0}(1785,2250)(1857,2250){1}
wire w441;    //: /sn:0 {0}(-414,764)(-414,803)(-242,803)(43:-242,828){1}
wire w796;    //: /sn:0 {0}(-551,1487)(-551,1470)(-520,1470)(-520,1501)(-504,1501){1}
wire w1376;    //: /sn:0 {0}(1979,2436)(2033,2436){1}
wire w621;    //: /sn:0 {0}(1229,1222)(1289,1222){1}
wire w1459;    //: /sn:0 {0}(3341,2550)(3270,2550){1}
wire w123;    //: /sn:0 {0}(-281,330)(-281,262){1}
wire w56;    //: /sn:0 {0}(-873,366)(-935,366){1}
wire w691;    //: /sn:0 {0}(1857,1348)(1785,1348){1}
wire w359;    //: /sn:0 {0}(-1057,695)(-1117,695){1}
wire w1413;    //: /sn:0 {0}(882,2439)(936,2439){1}
wire Cr5;    //: /sn:0 {0}(1229,561)(3939,561)(3939,2452)(4095,2452){1}
wire w1417;    //: /sn:0 {0}(974,2517)(974,2476){1}
wire w408;    //: /sn:0 {0}(1058,893)(1107,893){1}
wire w1220;    //: /sn:0 {0}(622,2069)(622,2023){1}
wire w1024;    //: /sn:0 {0}(1663,1800)(1591,1800){1}
wire w381;    //: /sn:0 {0}(143,601)(143,639)(310,639)(43:310,659){1}
wire A8;    //: {0}(3:2069,1315)(2069,-81)(1082,-81)(1082,-293){1}
wire w1498;    //: /sn:0 {0}(1701,2517)(1701,2476){1}
wire w1291;    //: /sn:0 {0}(2490,2322)(2490,2354)(2668,2354)(24:2668,2371){1}
wire w941;    //: /sn:0 {0}(-135,1650)(-197,1650){1}
wire w340;    //: /sn:0 {0}(-567,727)(-504,727){1}
wire w1328;    //: /sn:0 {0}(539,2285)(584,2285){1}
wire w269;    //: /sn:0 {0}(-1421,532)(-1483,532){1}
wire w54;    //: /sn:0 {0}(355,363)(417,363){1}
wire w647;    //: /sn:0 {0}(-504,1193)(-567,1193){1}
wire w1281;    //: /sn:0 {0}(2033,2250)(1979,2250){1}
wire w884;    //: /sn:0 {0}(2303,1719)(2303,1751)(2473,1751)(30:2473,1767){1}
wire w1067;    //: /sn:0 {0}(1229,1951)(1289,1951){1}
wire w110;    //: /sn:0 {0}(147,262)(147,311)(310,311)(24:310,330){1}
wire w46;    //: /sn:0 {0}(760,363)(706,363){1}
wire w532;    //: /sn:0 {0}(-197,1066)(-135,1066){1}
wire w968;    //: /sn:0 {0}(853,1719)(853,1749)(1013,1749)(30:1013,1767){1}
wire w1461;    //: /sn:0 {0}(4100,2693)(3379,2693)(3379,2622){1}
wire w787;    //: /sn:0 {0}(2033,1500)(1979,1500){1}
wire w1493;    //: /sn:0 {0}(30:1934,2517)(1934,2502)(1756,2502)(1756,2476){1}
wire w136;    //: /sn:0 {0}(-1933,262)(-1933,277){1}
wire w893;    //: /sn:0 {0}(-365,1698)(-365,1718)(-336,1718)(-336,1682)(-319,1682){1}
wire w1529;    //: /sn:0 {0}(24:1366,2517)(1366,2504)(1201,2504)(1201,2476){1}
wire w1009;    //: /sn:0 {0}(539,1801)(585,1801){1}
wire w357;    //: /sn:0 {0}(-1117,727)(-1057,727){1}
wire w735;    //: /sn:0 {0}(1058,1380)(1107,1380){1}
wire w1483;    //: /sn:0 {0}(2874,2622)(2874,2634){1}
wire w832;    //: /sn:0 {0}(1289,1500)(1229,1500){1}
wire A7;    //: {0}(3:2246,1467)(2246,-103)(1101,-103)(1101,-293){1}
wire w83;    //: /sn:0 {0}(760,529)(706,529){1}
wire w839;    //: /sn:0 {0}(-135,1503)(-197,1503){1}
wire w1455;    //: /sn:0 {0}(2033,2582)(1979,2582){1}
wire w918;    //: /sn:0 {0}(-25:974,1614)(974,1572){1}
wire w309;    //: /sn:0 {0}(1145,828)(1145,764){1}
wire w492;    //: /sn:0 {0}(53,1031)(-13,1031){1}
wire w26;    //: /sn:0 {0}(-689,222)(-751,222){1}
wire w1164;    //: /sn:0 {0}(1289,2102)(1229,2102){1}
wire w13;    //: /sn:0 {0}(-967,262)(-967,309)(-796,309)(43:-796,330){1}
wire w321;    //: /sn:0 {0}(233,692)(175,692){1}
wire w1467;    //: /sn:0 {0}(4100,2703)(3186,2703)(3186,2622){1}
wire w1381;    //: /sn:0 {0}(2155,2436)(2210,2436){1}
wire w1131;    //: /sn:0 {0}(62:130,1918)(130,1900)(-47,1900)(-47,1872){1}
wire w59;    //: /sn:0 {0}(-1019,435)(-25:-1019,496){1}
wire w25;    //: /sn:0 {0}(622,330)(622,262){1}
wire w423;    //: /sn:0 {0}(-25:798,828)(798,764){1}
wire w765;    //: /sn:0 {0}(43:1013,1315)(1013,1293)(850,1293)(850,1262){1}
wire w901;    //: /sn:0 {0}(1229,1679)(1289,1679){1}
wire w498;    //: /sn:0 {0}(1411,1063)(1469,1063){1}
wire w1162;    //: /sn:0 {0}(1229,2134)(1289,2134){1}
wire w36;    //: /sn:0 {0}(-25:-1201,330)(-1201,262){1}
wire w60;    //: /sn:0 {0}(-935,398)(-873,398){1}
wire w1068;    //: /sn:0 {0}(1107,1951)(1058,1951){1}
wire w949;    //: /sn:0 {0}(62:1934,1614)(1934,1596)(1751,1596)(1751,1572){1}
wire w1108;    //: /sn:0 {0}(882,1986)(936,1986){1}
wire w608;    //: /sn:0 {0}(539,1222)(584,1222){1}
wire w996;    //: /sn:0 {0}(-25:1327,1918)(1327,1872){1}
wire w179;    //: /sn:0 {0}(-13,395)(53,395){1}
wire w1526;    //: /sn:0 {0}(3002,2517)(3002,2476){1}
wire w1481;    //: /sn:0 {0}(2902,2550)(2964,2550){1}
wire w1061;    //: /sn:0 {0}(2713,1951)(2780,1951){1}
wire w421;    //: /sn:0 {0}(355,893)(417,893){1}
wire w1;    //: /sn:0 {0}(321,262)(321,309)(494,309)(62:494,330){1}
wire w396;    //: /sn:0 {0}(-135,861)(-197,861){1}
wire w194;    //: /sn:0 {0}(-1699,435)(-1699,468)(-1528,468)(62:-1528,496){1}
wire w912;    //: /sn:0 {0}(584,1650)(539,1650){1}
wire w874;    //: /sn:0 {0}(706,1679)(760,1679){1}
wire w504;    //: /sn:0 {0}(1229,1063)(1289,1063){1}
wire w1186;    //: /sn:0 {0}(1591,2102)(1663,2102){1}
wire w27;    //: /sn:0 {0}(-651,330)(-651,262){1}
wire w687;    //: /sn:0 {0}(584,1380)(539,1380){1}
wire w80;    //: /sn:0 {0}(2332,1532)(3845,1532)(3845,2512)(4095,2512){1}
wire w965;    //: /sn:0 {0}(2518,1800)(2591,1800){1}
wire w646;    //: /sn:0 {0}(-382,1193)(-319,1193){1}
wire w1341;    //: /sn:0 {0}(43:2110,2217)(2110,2201)(1947,2201)(1947,2174){1}
wire w415;    //: /sn:0 {0}(271,764)(271,828){1}
wire w544;    //: /sn:0 {0}(760,1031)(706,1031){1}
wire w971;    //: /sn:0 {0}(1058,1800)(1107,1800){1}
wire w1023;    //: /sn:0 {0}(1591,1832)(1663,1832){1}
wire w425;    //: /sn:0 {0}(882,861)(936,861){1}
wire w512;    //: /sn:0 {0}(355,1063)(417,1063){1}
wire w591;    //: /sn:0 {0}(417,1222)(355,1222){1}
wire w1176;    //: /sn:0 {0}(2518,2134)(2591,2134){1}
wire w465;    //: /sn:0 {0}(-1149,764)(-1149,804)(-980,804)(43:-980,828){1}
wire w350;    //: /sn:0 {0}(455,601)(455,659){1}
wire w1197;    //: /sn:0 {0}(2332,2134)(2396,2134){1}
wire w1471;    //: /sn:0 {0}(2248,2517)(2248,2476){1}
wire w1349;    //: /sn:0 {0}(3270,2404)(3341,2404){1}
wire w133;    //: /sn:0 {0}(-1787,193)(-1816,193)(-1816,193)(-1849,193){1}
wire w1008;    //: /sn:0 {0}(760,1803)(706,1803){1}
wire w513;    //: /sn:0 {0}(584,1031)(539,1031){1}
wire Cr8;    //: /sn:0 {0}(-935,564)(-873,564){1}
wire w705;    //: /sn:0 {0}(936,1348)(882,1348){1}
wire w1503;    //: /sn:0 {0}(2518,2582)(2591,2582){1}
wire w229;    //: /sn:0 {0}(-13,561)(53,561){1}
wire w303;    //: /sn:0 {0}(-135,724)(-197,724){1}
wire w585;    //: /sn:0 {0}(271,1103)(271,1157){1}
wire w128;    //: /sn:0 {0}(-416,262)(-416,309)(-242,309)(62:-242,330){1}
wire w682;    //: /sn:0 {0}(355,1380)(417,1380){1}
wire w188;    //: /sn:0 {0}(-1328,435)(-1328,472)(-1162,472)(30:-1162,496){1}
wire w533;    //: /sn:0 {0}(147,933)(147,972)(310,972)(24:310,998){1}
wire w1216;    //: /sn:0 {0}(2033,2102)(1979,2102){1}
wire w1193;    //: /sn:0 {0}(2332,2102)(2396,2102){1}
wire w464;    //: /sn:0 {0}(-1117,896)(-1057,896){1}
wire w185;    //: /sn:0 {0}(-1483,398)(-1421,398){1}
wire w195;    //: /sn:0 {0}(-1749,435)(-1749,450){1}
wire w644;    //: /sn:0 {0}(-466,1103)(-466,1157){1}
wire Cr30;    //: /sn:0 {0}(1058,2285)(1107,2285){1}
wire w908;    //: /sn:0 {0}(1701,1767)(1701,1719){1}
wire w1265;    //: /sn:0 {0}(3002,2217)(3002,2174){1}
wire w791;    //: /sn:0 {0}(1895,1467)(1895,1420){1}
wire Cr31;    //: /sn:0 {0}(3650,2582)(4095,2582){1}
wire w1502;    //: /sn:0 {0}(2629,2517)(2629,2476){1}
wire w86;    //: /sn:0 {0}(2713,1832)(3824,1832)(3824,2532)(4095,2532){1}
wire w349;    //: /sn:0 {0}(326,601)(326,638)(494,638)(30:494,659){1}
wire w1489;    //: /sn:0 {0}(1411,2551)(1469,2551){1}
wire w1439;    //: /sn:0 {0}(43:2473,2517)(2473,2501)(2300,2501)(2300,2476){1}
wire w742;    //: /sn:0 {0}(-197,1351)(-135,1351){1}
wire Cr22;    //: /sn:0 {0}(355,1682)(417,1682){1}
wire w1325;    //: /sn:0 {0}(584,2253)(539,2253){1}
wire w1531;    //: /sn:0 {0}(1383,2622)(1383,2634){1}
wire w1063;    //: /sn:0 {0}(2818,2069)(2818,2023){1}
wire w8;    //: /sn:0 {0}(507,262)(507,309)(661,309)(43:661,330){1}
wire w140;    //: /sn:0 {0}(-1421,225)(-1443,225)(-1443,225)(-1483,225){1}
wire w147;    //: /sn:0 {0}(-1605,193)(-1629,193)(-1629,193)(-1665,193){1}
wire w1201;    //: /sn:0 {0}(882,2103)(936,2103){1}
wire w44;    //: /sn:0 {0}(-504,395)(-567,395){1}
wire w604;    //: /sn:0 {0}(-928,1175)(-928,1158)(-890,1158)(-890,1191)(-873,1191){1}
wire w659;    //: /sn:0 {0}(43:-427,1315)(-427,1293)(-599,1293)(-599,1262){1}
wire w797;    //: /sn:0 {0}(-549,1551)(-549,1571)(-520,1571)(-520,1535)(-504,1535){1}
wire w1081;    //: /sn:0 {0}(2396,1951)(2332,1951){1}
wire w14;    //: /sn:0 {0}(-1299,191)(-1253,191)(-1253,191)(-1239,191){1}
wire w45;    //: /sn:0 {0}(706,395)(760,395){1}
wire w1495;    //: /sn:0 {0}(2127,2622)(2127,2634){1}
wire w1260;    //: /sn:0 {0}(1469,2250)(1411,2250){1}
wire w74;    //: /sn:0 {0}(-504,529)(-567,529){1}
wire w1097;    //: /sn:0 {0}(2155,1951)(2210,1951){1}
wire w129;    //: /sn:0 {0}(-25:-466,330)(-466,262){1}
wire w610;    //: /sn:0 {0}(539,1190)(584,1190){1}
wire A1;    //: {0}(1:3377,2371)(3377,-240)(1237,-240)(1237,-293){1}
wire w1200;    //: /sn:0 {0}(1107,2105)(1058,2105){1}
wire w675;    //: /sn:0 {0}(2033,1380)(1979,1380){1}
wire w1350;    //: /sn:0 {0}(3435,2476)(3435,2495)(3605,2495)(24:3605,2517){1}
wire w15;    //: /sn:0 {0}(539,222)(584,222){1}
wire w994;    //: /sn:0 {0}(1229,1800)(1289,1800){1}
wire w455;    //: /sn:0 {0}(-873,864)(-935,864){1}
wire w792;    //: /sn:0 {0}(1785,1532)(1857,1532){1}
wire w1532;    //: /sn:0 {0}(4100,2803)(1327,2803)(1327,2622){1}
wire w934;    //: /sn:0 {0}(175,1650)(233,1650){1}
wire w989;    //: /sn:0 {0}(-188,1851)(-188,1872)(-156,1872)(-156,1835)(-135,1835){1}
wire A0;    //: {0}(1:3564,2517)(3564,-264)(1258,-264)(1258,-293){1}
wire w1090;    //: /sn:0 {0}(1411,1951)(1469,1951){1}
wire w307;    //: /sn:0 {0}(1107,692)(1058,692){1}
wire w749;    //: /sn:0 {0}(-504,1351)(-567,1351){1}
wire w836;    //: /sn:0 {0}(-97,1420)(-97,1467){1}
wire w306;    //: /sn:0 {0}(1058,724)(1107,724){1}
wire w755;    //: /sn:0 {0}(-414,1420)(-414,1449)(-242,1449)(43:-242,1467){1}
wire w1268;    //: /sn:0 {0}(3057,2322)(3057,2352)(3225,2352)(30:3225,2371){1}
wire w458;    //: /sn:0 {0}(-689,896)(-751,896){1}
wire w810;    //: /sn:0 {0}(1411,1500)(1469,1500){1}
wire w418;    //: /sn:0 {0}(175,861)(233,861){1}
wire w299;    //: /sn:0 {0}(-197,692)(-135,692){1}
wire B13;    //: {0}(20:-1528,157)(-1528,-238)(534,-238)(534,-294){1}
wire w793;    //: /sn:0 {0}(1857,1500)(1785,1500){1}
wire w640;    //: /sn:0 {0}(936,1190)(882,1190){1}
wire w875;    //: /sn:0 {0}(882,1647)(936,1647){1}
wire A13;    //: {0}(13:1143,496)(1143,47)(990,47)(990,-293){1}
wire w1446;    //: /sn:0 {0}(3622,2622)(3622,2634){1}
wire w548;    //: /sn:0 {0}(-651,933)(-651,998){1}
wire w601;    //: /sn:0 {0}(1469,1190)(1411,1190){1}
wire w944;    //: /sn:0 {0}(-197,1682)(-135,1682){1}
wire w1052;    //: /sn:0 {0}(455,1918)(455,1872){1}
wire w369;    //: /sn:0 {0}(-1331,601)(-1331,643)(-1162,643)(43:-1162,659){1}
wire w66;    //: /sn:0 {0}(-25:455,496)(455,435){1}
wire w73;    //: /sn:0 {0}(-382,529)(-319,529){1}
wire w1519;    //: /sn:0 {0}(4100,2833)(795,2833)(795,2622){1}
wire w609;    //: /sn:0 {0}(760,1190)(706,1190){1}
wire w656;    //: /sn:0 {0}(-751,1225)(-689,1225){1}
wire w813;    //: /sn:0 {0}(1593,1532)(1663,1532){1}
wire w1302;    //: /sn:0 {0}(-25:1701,2217)(1701,2174){1}
wire w938;    //: /sn:0 {0}(233,1682)(175,1682){1}
wire w1499;    //: /sn:0 {0}(1753,2622)(1753,2632){1}
wire w285;    //: /sn:0 {0}(-45,435)(-45,472)(130,472)(43:130,496){1}
wire w256;    //: /sn:0 {0}(233,529)(175,529){1}
wire w1085;    //: /sn:0 {0}(-4,2000)(-4,2019)(32,2019)(32,1986)(53,1986){1}
wire w1064;    //: /sn:0 {0}(30:1184,1918)(1184,1902)(1029,1902)(1029,1872){1}
wire B12;    //: {0}(20:-1344,157)(-1344,-223)(561,-223)(561,-294){1}
wire w1079;    //: /sn:0 {0}(2434,1872)(2434,1918){1}
wire w988;    //: /sn:0 {0}(-190,1787)(-190,1770)(-157,1770)(-157,1801)(-135,1801){1}
wire w709;    //: /sn:0 {0}(882,1380)(936,1380){1}
wire w466;    //: /sn:0 {0}(-1019,764)(-1019,828){1}
wire w906;    //: /sn:0 {0}(1591,1647)(1663,1647){1}
wire w1277;    //: /sn:0 {0}(370,2299)(370,2319)(398,2319)(398,2285)(417,2285){1}
wire w477;    //: /sn:0 {0}(323,764)(323,806)(494,806)(43:494,828){1}
wire w1001;    //: /sn:0 {0}(1979,1800)(2033,1800){1}
wire w33;    //: /sn:0 {0}(936,395)(882,395){1}
wire w453;    //: /sn:0 {0}(-935,896)(-873,896){1}
wire w1157;    //: /sn:0 {0}(2902,2102)(2964,2102){1}
wire w490;    //: /sn:0 {0}(-13,1063)(53,1063){1}
wire w126;    //: /sn:0 {0}(-567,222)(-507,222)(-507,222)(-504,222){1}
wire w365;    //: /sn:0 {0}(-1239,695)(-1299,695){1}
wire w509;    //: /sn:0 {0}(-1124,1082)(-1124,1102)(-1085,1102)(-1085,1066)(-1057,1066){1}
wire w963;    //: /sn:0 {0}(2591,1832)(2518,1832){1}
wire w220;    //: /sn:0 {0}(-1678,515)(-1678,498)(-1633,498)(-1633,530)(-1605,530){1}
wire w79;    //: /sn:0 {0}(936,529)(882,529){1}
wire w1051;    //: /sn:0 {0}(24:661,1918)(661,1901)(511,1901)(511,1872){1}
wire w529;    //: /sn:0 {0}(-382,1032)(-319,1032){1}
wire w882;    //: /sn:0 {0}(2155,1679)(2210,1679){1}
wire w1418;    //: /sn:0 {0}(1107,2439)(1058,2439){1}
wire w998;    //: /sn:0 {0}(1757,1719)(1757,1750)(1934,1750)(24:1934,1767){1}
wire w993;    //: /sn:0 {0}(1469,1800)(1411,1800){1}
wire w837;    //: /sn:0 {0}(-197,1535)(-135,1535){1}
wire w1084;    //: /sn:0 {0}(-6,1936)(-6,1918)(32,1918)(32,1952)(53,1952){1}
wire A3;    //: {0}(1:3000,2069)(3000,-196)(1186,-196)(1186,-293){1}
wire w1092;    //: /sn:0 {0}(-25:1507,2069)(1507,2023){1}
wire w1490;    //: /sn:0 {0}(1557,2622)(1557,2631){1}
wire w1139;    //: /sn:0 {0}(323,2023)(323,2050)(494,2050)(43:494,2069){1}
wire w387;    //: /sn:0 {0}(1469,893)(1411,893){1}
wire w109;    //: /sn:0 {0}(-13,190)(53,190){1}
wire w164;    //: /sn:0 {0}(-197,395)(-135,395){1}
wire w223;    //: /sn:0 {0}(-97,435)(-97,496){1}
wire w237;    //: /sn:0 {0}(539,561)(584,561){1}
wire w560;    //: /sn:0 {0}(-935,1066)(-873,1066){1}
wire w820;    //: /sn:0 {0}(355,1535)(417,1535){1}
wire w325;    //: /sn:0 {0}(175,724)(233,724){1}
wire w616;    //: /sn:0 {0}(1107,1222)(1058,1222){1}
wire w658;    //: /sn:0 {0}(-651,1103)(-651,1157){1}
wire w842;    //: /sn:0 {0}(53,1535)(-13,1535){1}
wire B14;    //: {0}(19:-1710,157)(-1710,-254)(507,-254)(507,-294){1}
wire w1465;    //: /sn:0 {0}(3148,2550)(3086,2550){1}
wire w624;    //: /sn:0 {0}(53,1193)(-13,1193){1}
wire A10;    //: {0}(6:1699,998)(1699,-39)(1047,-39)(1047,-293){1}
wire w1293;    //: /sn:0 {0}(2518,2282)(2591,2282){1}
wire w180;    //: /sn:0 {0}(53,363)(-13,363){1}
wire w1368;    //: /sn:0 {0}(2902,2436)(2964,2436){1}
wire B1;    //: {0}(59:661,157)(661,48)(819,48)(819,-294){1}
wire w1500;    //: /sn:0 {0}(4100,2783)(1701,2783)(1701,2622){1}
wire w1213;    //: /sn:0 {0}(1950,2023)(1950,2051)(2110,2051)(30:2110,2069){1}
wire w979;    //: /sn:0 {0}(2396,1800)(2332,1800){1}
wire w1088;    //: /sn:0 {0}(1411,1983)(1469,1983){1}
wire w233;    //: /sn:0 {0}(539,529)(584,529){1}
wire w1125;    //: /sn:0 {0}(355,1986)(417,1986){1}
wire w35;    //: /sn:0 {0}(-1151,262)(-1151,306)(-980,306)(62:-980,330){1}
wire w153;    //: /sn:0 {0}(-1697,262)(-1697,298)(-1528,298)(43:-1528,330){1}
wire w867;    //: /sn:0 {0}(2396,1679)(2332,1679){1}
wire Cr16;    //: /sn:0 {0}(-197,1225)(-135,1225){1}
wire w1359;    //: /sn:0 {0}(1857,2436)(1785,2436){1}
wire w1232;    //: /sn:0 {0}(355,2137)(417,2137){1}
wire w771;    //: /sn:0 {0}(2210,1532)(2155,1532){1}
wire w1000;    //: /sn:0 {0}(1857,1832)(1785,1832){1}
wire w127;    //: /sn:0 {0}(-567,190)(-507,190)(-507,190)(-504,190){1}
wire w416;    //: /sn:0 {0}(175,893)(233,893){1}
wire w55;    //: /sn:0 {0}(355,395)(417,395){1}
wire w645;    //: /sn:0 {0}(-567,1225)(-504,1225){1}
wire w1130;    //: /sn:0 {0}(584,1986)(539,1986){1}
wire w1506;    //: /sn:0 {0}(4100,2733)(2629,2733)(2629,2622){1}
wire w1327;    //: /sn:0 {0}(455,2322)(455,2337){1}
wire w1076;    //: /sn:0 {0}(2684,2023)(2684,2055)(2857,2055)(30:2857,2069){1}
wire w114;    //: /sn:0 {0}(-197,222)(-133,222)(-133,222)(-135,222){1}
wire w1222;    //: /sn:0 {0}(706,2105)(760,2105){1}
wire w143;    //: /sn:0 {0}(-1383,262)(-1383,330){1}
wire w869;    //: /sn:0 {0}(2332,1647)(2396,1647){1}
wire w1177;    //: /sn:0 {0}(2591,2102)(2518,2102){1}
wire w888;    //: /sn:0 {0}(1979,1679)(2033,1679){1}
wire w1475;    //: /sn:0 {0}(2298,2622)(2298,2631){1}
wire w1453;    //: /sn:0 {0}(1950,2622)(1950,2632){1}
wire Cr18;    //: /sn:0 {0}(-13,1383)(53,1383){1}
wire w1363;    //: /sn:0 {0}(3148,2404)(3086,2404){1}
wire w1259;    //: /sn:0 {0}(1591,2250)(1663,2250){1}
wire w1258;    //: /sn:0 {0}(1411,2282)(1469,2282){1}
wire w1089;    //: /sn:0 {0}(1663,1951)(1591,1951){1}
wire w1285;    //: /sn:0 {0}(1979,2282)(2033,2282){1}
wire w1066;    //: /sn:0 {0}(1058,1983)(1107,1983){1}
wire w978;    //: /sn:0 {0}(2332,1832)(2396,1832){1}
wire w1311;    //: /sn:0 {0}(2155,2282)(2210,2282){1}
wire w367;    //: /sn:0 {0}(-1383,764)(-1383,779){1}
wire w206;    //: /sn:0 {0}(-1201,435)(-1201,496){1}
wire w520;    //: /sn:0 {0}(936,1063)(882,1063){1}
wire w10;    //: /sn:0 {0}(-1117,225)(-1063,225)(-1063,225)(-1057,225){1}
wire w111;    //: /sn:0 {0}(91,330)(91,262){1}
wire w1127;    //: /sn:0 {0}(417,1954)(355,1954){1}
wire w436;    //: /sn:0 {0}(-382,896)(-319,896){1}
wire w514;    //: /sn:0 {0}(355,1031)(417,1031){1}
wire w697;    //: /sn:0 {0}(1663,1348)(1591,1348){1}
wire w904;    //: /sn:0 {0}(1663,1679)(1591,1679){1}
wire w389;    //: /sn:0 {0}(1411,861)(1469,861){1}
wire w1384;    //: /sn:0 {0}(2591,2436)(2518,2436){1}
wire w1080;    //: /sn:0 {0}(2332,1983)(2396,1983){1}
wire w970;    //: /sn:0 {0}(882,1832)(936,1832){1}
wire w200;    //: /sn:0 {0}(-1567,496)(-1567,435){1}
wire w1012;    //: /sn:0 {0}(706,1835)(760,1835){1}
wire w17;    //: /sn:0 {0}(677,262)(677,310)(837,310)(30:837,330){1}
wire w1215;    //: /sn:0 {0}(1979,2134)(2033,2134){1}
wire w1192;    //: /sn:0 {0}(2210,2134)(2155,2134){1}
wire w49;    //: /sn:0 {0}(539,395)(584,395){1}
wire w706;    //: /sn:0 {0}(706,1348)(760,1348){1}
wire w1450;    //: /sn:0 {0}(1785,2582)(1857,2582){1}
wire w1472;    //: /sn:0 {0}(2155,2582)(2210,2582){1}
wire w587;    //: /sn:0 {0}(355,1190)(417,1190){1}
wire Cr26;    //: /sn:0 {0}(706,1986)(760,1986){1}
wire w160;    //: /sn:0 {0}(-135,363)(-197,363){1}
wire w64;    //: /sn:0 {0}(-835,435)(-835,496){1}
wire w362;    //: /sn:0 {0}(-873,727)(-935,727){1}
wire w312;    //: /sn:0 {0}(882,724)(936,724){1}
wire w298;    //: /sn:0 {0}(-382,724)(-319,724){1}
wire w271;    //: /sn:0 {0}(-1567,601)(-1567,616){1}
//: enddecls

  HD g8 (.B(B9), .A(w1444), .CrIn(w22), .PrIn(w21), .PrOut(w12), .BOut(w30), .Q(w31), .CrOut(w26));   //: @(-872, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>111 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g164 (.B(w825), .A(w686), .CrIn(w820), .PrIn(w780), .PrOut(w816), .BOut(w827), .Q(w911), .CrOut(w778));   //: @(418, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  assign A9 = A[9]; //: TAP g312 @(1064,-299) /sn:0 /R:1 /w:[ 1 20 19 ] /ss:1
  HD g258 (.B(w1235), .A(w1225), .CrIn(w1328), .PrIn(w1319), .PrOut(w1325), .BOut(w1331), .Q(w1420), .CrOut(w1317));   //: @(585, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g224 (.B(w1141), .A(w987), .CrIn(w1101), .PrIn(w1081), .PrOut(w1097), .BOut(w1237), .Q(w1191), .CrOut(w1080));   //: @(2211, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g226 (.B(w1055), .A(w1150), .CrIn(w1093), .PrIn(w1120), .PrOut(w1089), .BOut(w1245), .Q(w1152), .CrOut(w1119));   //: @(1664, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g243 (.B(w1147), .A(w1242), .CrIn(w1226), .PrIn(w1201), .PrOut(w1222), .BOut(w1243), .Q(w1244), .CrOut(Cr28));   //: @(761, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  assign B3 = B[3]; //: TAP g30 @(775,-300) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  HD g92 (.B(w441), .A(w442), .CrIn(w436), .PrIn(w396), .PrOut(w432), .BOut(w443), .Q(w527), .CrOut(w394));   //: @(-318, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g74 (.B(w345), .A(w346), .CrIn(w340), .PrIn(w300), .PrOut(w336), .BOut(w441), .Q(w348), .CrOut(w298));   //: @(-503, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g198 (.B(w1006), .A(w924), .CrIn(Cr24), .PrIn(w1008), .PrOut(w1009), .BOut(w1010), .Q(w1011), .CrOut(w1012));   //: @(586, 1768) /sz:(119, 104) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  NandNOT g1 (.in1(w4), .out(w104));   //: @(-2072, 177) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g130 (.B(w552), .A(w644), .CrIn(w645), .PrIn(w646), .PrOut(w647), .BOut(w648), .Q(w649), .CrOut(w650));   //: @(-503, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g183 (.B(w925), .A(w926), .CrIn(w927), .PrIn(w906), .PrOut(w928), .BOut(w1021), .Q(w1054), .CrOut(w904));   //: @(1470, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g111 (.B(w449), .A(w428), .CrIn(w543), .PrIn(w522), .PrOut(w544), .BOut(w545), .Q(w670), .CrOut(w520));   //: @(761, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g253 (.B(w1207), .A(w1302), .CrIn(w1263), .PrIn(w1282), .PrOut(w1259), .BOut(w1397), .Q(w1304), .CrOut(w1280));   //: @(1664, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g274 (.B(w1320), .A(w1412), .CrIn(w1413), .PrIn(w1414), .PrOut(w1415), .BOut(w1507), .Q(w1417), .CrOut(w1418));   //: @(937, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g260 (.B(w1239), .A(w1334), .CrIn(w1293), .PrIn(w1273), .PrOut(w1289), .BOut(w1335), .Q(w1383), .CrOut(w1272));   //: @(2592, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g179 (.B(w811), .A(w856), .CrIn(w904), .PrIn(w905), .PrOut(w906), .BOut(w998), .Q(w908), .CrOut(w909));   //: @(1664, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g70 (.B(w227), .A(w288), .CrIn(w320), .PrIn(w321), .PrOut(w322), .BOut(w323), .Q(w438), .CrOut(w325));   //: @(54, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g206 (.B(w1045), .A(w891), .CrIn(w1005), .PrIn(w985), .PrOut(w1001), .BOut(w1141), .Q(w1095), .CrOut(w984));   //: @(2034, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g10 (.B(B11), .A(w1444), .CrIn(Cr6), .PrIn(w6), .PrOut(w14), .BOut(w35), .Q(w36), .CrOut(w10));   //: @(-1238, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>115 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g25 (.B(B4), .A(w1444), .CrIn(w107), .PrIn(w9), .PrOut(w109), .BOut(w110), .Q(w111), .CrOut(w2));   //: @(54, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>101 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g149 (.B(w654), .A(w748), .CrIn(w701), .PrIn(w749), .PrOut(w700), .BOut(w843), .Q(w751), .CrOut(w752));   //: @(-688, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g64 (.B(w285), .A(w286), .CrIn(w229), .PrIn(w256), .PrOut(w225), .BOut(w381), .Q(w288), .CrOut(w255));   //: @(54, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g220 (.B(w1032), .A(w1052), .CrIn(w1125), .PrIn(w1126), .PrOut(w1127), .BOut(w1128), .Q(w1129), .CrOut(w1130));   //: @(418, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g49 (.B(w142), .A(w36), .CrIn(w190), .PrIn(w57), .PrOut(w186), .BOut(w205), .Q(w206), .CrOut(Cr7));   //: @(-1238, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g270 (.B(w1390), .A(w1391), .CrIn(Cr32), .PrIn(w1392), .PrOut(w1393), .BOut(w1486), .Q(w1530), .CrOut(w1396));   //: @(1290, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  assign A12 = A[12]; //: TAP g35 @(1008,-299) /sn:0 /R:1 /w:[ 1 26 25 ] /ss:1
  HD g181 (.B(w917), .A(w918), .CrIn(w879), .PrIn(w898), .PrOut(w875), .BOut(w919), .Q(w920), .CrOut(w896));   //: @(937, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g85 (.B(w400), .A(w308), .CrIn(w402), .PrIn(w389), .PrOut(w403), .BOut(w496), .Q(w503), .CrOut(w387));   //: @(1290, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g67 (.B(w304), .A(w71), .CrIn(w306), .PrIn(w293), .PrOut(w307), .BOut(w400), .Q(w309), .CrOut(w291));   //: @(1108, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g192 (.B(w968), .A(w920), .CrIn(w970), .PrIn(w971), .PrOut(w972), .BOut(w1064), .Q(w974), .CrOut(w975));   //: @(937, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g126 (.B(w622), .A(w623), .CrIn(Cr16), .PrIn(w624), .PrOut(w625), .BOut(w718), .Q(w762), .CrOut(w628));   //: @(-134, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  assign A14 = A[14]; //: TAP g33 @(972,-299) /sn:0 /R:1 /w:[ 1 30 29 ] /ss:1
  assign B6 = B[6]; //: TAP g300 @(712,-300) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  HD g54 (.B(w58), .A(w64), .CrIn(Cr8), .PrIn(w240), .PrOut(w241), .BOut(w242), .Q(w378), .CrOut(w244));   //: @(-872, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g234 (.B(w1106), .A(w1199), .CrIn(Cr28), .PrIn(w1200), .PrOut(w1201), .BOut(w1202), .Q(w1338), .CrOut(w1204));   //: @(937, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g132 (.B(w563), .A(w658), .CrIn(w656), .PrIn(w647), .PrOut(w653), .BOut(w659), .Q(w748), .CrOut(w645));   //: @(-688, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g163 (.B(w821), .A(w822), .CrIn(w783), .PrIn(w802), .PrOut(w779), .BOut(w917), .Q(w873), .CrOut(w800));   //: @(761, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g12 (.B(w30), .A(w27), .CrIn(w39), .PrIn(w40), .PrOut(w41), .BOut(w42), .Q(w43), .CrOut(w44));   //: @(-688, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g217 (.B(w1109), .A(w996), .CrIn(w1071), .PrIn(w1090), .PrOut(w1067), .BOut(w1111), .Q(w1161), .CrOut(w1088));   //: @(1290, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g222 (.B(w1043), .A(w1033), .CrIn(w1136), .PrIn(w1127), .PrOut(w1133), .BOut(w1139), .Q(w1228), .CrOut(w1125));   //: @(234, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g298 (.B(w1439), .A(w1410), .CrIn(w1477), .PrIn(w1504), .PrOut(w1473), .BOut(w1535), .Q(w1536), .CrOut(w1503));   //: @(2397, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g106 (.B(w419), .A(w480), .CrIn(w512), .PrIn(w513), .PrOut(w514), .BOut(w515), .Q(w630), .CrOut(w517));   //: @(418, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  NandNOT g177 (.in1(w892), .out(w893));   //: @(-389, 1635) /sz:(46, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g194 (.B(w982), .A(w885), .CrIn(w984), .PrIn(w979), .PrOut(w985), .BOut(w986), .Q(w987), .CrOut(w978));   //: @(2211, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g230 (.B(w1174), .A(w1175), .CrIn(w1176), .PrIn(w1171), .PrOut(w1177), .BOut(w1178), .Q(w1334), .CrOut(w1170));   //: @(2592, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  assign B13 = B[13]; //: TAP g307 @(534,-300) /sn:0 /R:1 /w:[ 1 28 27 ] /ss:1
  HD g228 (.B(w1069), .A(w1161), .CrIn(w1162), .PrIn(w1163), .PrOut(w1164), .BOut(w1165), .Q(w1166), .CrOut(w1167));   //: @(1290, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  //: joint g19 (w1444) @(1819, 1031) /w:[ 40 39 82 -1 ]
  HD g114 (.B(w561), .A(w457), .CrIn(w560), .PrIn(w551), .PrOut(w557), .BOut(w563), .Q(w652), .CrOut(w549));   //: @(-872, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g196 (.B(w899), .A(w991), .CrIn(w992), .PrIn(w993), .PrOut(w994), .BOut(w995), .Q(w996), .CrOut(w997));   //: @(1290, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  assign R = {w1519, w1524, w1513, w1532, w1491, w1500, w1454, w1496, w1476, w1536, w1506, w1484, w1528, w1467, w1461, w1447}; //: CONCAT g339  @(4105,2758) /sn:0 /w:[ 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  HD g125 (.B(w614), .A(w615), .CrIn(w616), .PrIn(w617), .PrOut(w618), .BOut(w710), .Q(w620), .CrOut(w621));   //: @(1108, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g281 (.B(w1350), .A(A0), .CrIn(w1443), .PrIn(w1444), .PrOut(w1445), .BOut(w1446), .Q(w1447), .CrOut(Cr31));   //: @(3529, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>63 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g100 (.B(w477), .A(w354), .CrIn(w421), .PrIn(w448), .PrOut(w417), .BOut(w573), .Q(w480), .CrOut(w447));   //: @(418, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g93 (.B(w445), .A(w332), .CrIn(w447), .PrIn(w426), .PrOut(w448), .BOut(w449), .Q(w574), .CrOut(w424));   //: @(585, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g63 (.B(w205), .A(w59), .CrIn(w266), .PrIn(w241), .PrOut(w262), .BOut(w377), .Q(w284), .CrOut(Cr8));   //: @(-1056, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g331 (w1444) @(-837, 129) /w:[ 12 -1 11 110 ]
  HD g262 (.B(w1341), .A(w1342), .CrIn(w1285), .PrIn(w1312), .PrOut(w1281), .BOut(w1437), .Q(w1375), .CrOut(w1311));   //: @(2034, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g101 (.B(w390), .A(A10), .CrIn(w483), .PrIn(w1444), .PrOut(w485), .BOut(w577), .Q(w487), .CrOut(Cr13));   //: @(1664, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>83 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g0 (.B(B3), .A(w1444), .CrIn(w2), .PrIn(w3), .PrOut(w9), .BOut(w1), .Q(w5), .CrOut(w7));   //: @(234, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>99 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g211 (.B(w1072), .A(w1073), .CrIn(w1074), .PrIn(w1061), .PrOut(w1075), .BOut(w1076), .Q(w1175), .CrOut(w1059));   //: @(2592, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g215 (.B(w1094), .A(w1095), .CrIn(w1096), .PrIn(w1097), .PrOut(w1098), .BOut(w1190), .Q(w1100), .CrOut(w1101));   //: @(2034, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g244 (.B(w1245), .A(w1122), .CrIn(w1189), .PrIn(w1216), .PrOut(w1185), .BOut(w1341), .Q(w1279), .CrOut(w1215));   //: @(1858, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g37 (.B(B6), .A(w1444), .CrIn(w120), .PrIn(w115), .PrOut(w121), .BOut(w122), .Q(w123), .CrOut(w114));   //: @(-318, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>105 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g120 (.B(w584), .A(w585), .CrIn(w586), .PrIn(w587), .PrOut(w588), .BOut(w680), .Q(w590), .CrOut(w591));   //: @(234, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g76 (.B(w355), .A(w284), .CrIn(w357), .PrIn(w358), .PrOut(w359), .BOut(w360), .Q(w466), .CrOut(w362));   //: @(-1056, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  NandNOT g267 (.in1(w1372), .out(w1373));   //: @(500, 2392) /sz:(48, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g75 (.B(w349), .A(w350), .CrIn(w351), .PrIn(w330), .PrOut(w352), .BOut(w445), .Q(w354), .CrOut(w328));   //: @(418, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g44 (.B(w110), .A(w5), .CrIn(w167), .PrIn(w54), .PrOut(w168), .BOut(w169), .Q(w170), .CrOut(w55));   //: @(234, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g152 (.B(w663), .A(w603), .CrIn(w717), .PrIn(w697), .PrOut(w713), .BOut(w853), .Q(w760), .CrOut(w696));   //: @(1470, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g47 (.B(w135), .A(w154), .CrIn(w156), .PrIn(w193), .PrOut(w53), .BOut(w194), .Q(w195), .CrOut(w196));   //: @(-1786, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g16 (.B(w35), .A(w32), .CrIn(Cr7), .PrIn(w56), .PrOut(w57), .BOut(w58), .Q(w59), .CrOut(w60));   //: @(-1056, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g3 (.B(B1), .A(w1444), .CrIn(w15), .PrIn(w19), .PrOut(w11), .BOut(w17), .Q(w25), .CrOut(w23));   //: @(585, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>95 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  NandNOT g159 (.in1(w796), .out(w797));   //: @(-574, 1488) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: IN g26 (B) @(864,-298) /sn:0 /R:2 /w:[ 0 ]
  HD g284 (.B(w1370), .A(w1365), .CrIn(w1464), .PrIn(w1459), .PrOut(w1465), .BOut(w1466), .Q(w1467), .CrOut(w1458));   //: @(3149, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g109 (.B(w533), .A(w534), .CrIn(w495), .PrIn(w514), .PrOut(w491), .BOut(w629), .Q(w585), .CrOut(w512));   //: @(234, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g143 (.B(w710), .A(w664), .CrIn(w712), .PrIn(w713), .PrOut(w714), .BOut(w806), .Q(w716), .CrOut(w717));   //: @(1290, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g334 (w1444) @(-1385, 129) /w:[ 6 -1 5 116 ]
  assign B8 = B[8]; //: TAP g302 @(665,-300) /sn:0 /R:1 /w:[ 1 18 17 ] /ss:1
  HD g158 (.B(w790), .A(w791), .CrIn(w792), .PrIn(w787), .PrOut(w793), .BOut(w794), .Q(w795), .CrOut(w786));   //: @(1858, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g23 (.B(w47), .A(w38), .CrIn(w78), .PrIn(w69), .PrOut(w79), .BOut(w304), .Q(w81), .CrOut(w67));   //: @(937, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  assign A5 = A[5]; //: TAP g316 @(1142,-299) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  assign B15 = B[15]; //: TAP g309 @(481,-300) /sn:0 /R:1 /w:[ 1 32 31 ] /ss:1
  HD g127 (.B(w629), .A(w630), .CrIn(w591), .PrIn(w610), .PrOut(w587), .BOut(w631), .Q(w681), .CrOut(w608));   //: @(418, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g104 (.B(w502), .A(w503), .CrIn(w504), .PrIn(w499), .PrOut(w505), .BOut(w506), .Q(w507), .CrOut(w498));   //: @(1290, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g86 (.B(w314), .A(w309), .CrIn(w408), .PrIn(w403), .PrOut(w409), .BOut(w502), .Q(w566), .CrOut(w402));   //: @(1108, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g24 (.B(w217), .A(w218), .CrIn(w82), .PrIn(w79), .PrOut(w83), .BOut(w84), .Q(w374), .CrOut(w78));   //: @(761, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g39 (.B(B7), .A(w1444), .CrIn(w126), .PrIn(w121), .PrOut(w127), .BOut(w128), .Q(w129), .CrOut(w120));   //: @(-503, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>107 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  assign A11 = A[11]; //: TAP g310 @(1027,-299) /sn:0 /R:1 /w:[ 1 24 23 ] /ss:1
  HD g289 (.B(w1399), .A(w1380), .CrIn(w1455), .PrIn(w1474), .PrOut(w1451), .BOut(w1495), .Q(w1496), .CrOut(w1472));   //: @(2034, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g121 (.B(w500), .A(w487), .CrIn(w594), .PrIn(w581), .PrOut(w595), .BOut(w596), .Q(w597), .CrOut(w579));   //: @(1664, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g110 (.B(w443), .A(w538), .CrIn(w532), .PrIn(w492), .PrOut(w528), .BOut(w539), .Q(w623), .CrOut(w490));   //: @(-134, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g60 (.B(w199), .A(w189), .CrIn(w272), .PrIn(w263), .PrOut(w269), .BOut(w369), .Q(w364), .CrOut(w261));   //: @(-1420, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g250 (.B(w1278), .A(w1279), .CrIn(w1280), .PrIn(w1281), .PrOut(w1282), .BOut(w1374), .Q(w1284), .CrOut(w1285));   //: @(1858, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: OUT g340 (R) @(4164,2758) /sn:0 /w:[ 0 ]
  HD g257 (.B(w1323), .A(w1236), .CrIn(w1277), .PrIn(w1325), .PrOut(w1276), .BOut(w1419), .Q(w1327), .CrOut(w1328));   //: @(418, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g82 (.B(w381), .A(w382), .CrIn(w325), .PrIn(w352), .PrOut(w321), .BOut(w477), .Q(w415), .CrOut(w351));   //: @(234, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g248 (.B(w1178), .A(w1173), .CrIn(w1272), .PrIn(w1267), .PrOut(w1273), .BOut(w1274), .Q(w1430), .CrOut(w1266));   //: @(2781, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g323 (w1444) @(620, 129) /w:[ 28 -1 27 94 ]
  assign B12 = B[12]; //: TAP g306 @(561,-300) /sn:0 /R:1 /w:[ 1 26 25 ] /ss:1
  HD g272 (.B(w1307), .A(w1262), .CrIn(w1396), .PrIn(w1356), .PrOut(w1392), .BOut(w1497), .Q(w1404), .CrOut(w1354));   //: @(1470, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g94 (.B(w360), .A(w452), .CrIn(w453), .PrIn(w454), .PrOut(w455), .BOut(w456), .Q(w457), .CrOut(w458));   //: @(-872, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g245 (.B(w1158), .A(A2), .CrIn(w1251), .PrIn(w1444), .PrOut(w1253), .BOut(w1254), .Q(w1361), .CrOut(w89));   //: @(3147, 2218) /sz:(122, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>67 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g107 (.B(w427), .A(w519), .CrIn(w520), .PrIn(w521), .PrOut(w522), .BOut(w614), .Q(w638), .CrOut(w525));   //: @(937, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g166 (.B(w744), .A(w836), .CrIn(w837), .PrIn(w838), .PrOut(w839), .BOut(w840), .Q(w841), .CrOut(w842));   //: @(-134, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g216 (.B(w1010), .A(w1020), .CrIn(Cr26), .PrIn(w1104), .PrOut(w1105), .BOut(w1106), .Q(w1242), .CrOut(w1108));   //: @(761, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  assign B7 = B[7]; //: TAP g301 @(688,-300) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  //: joint g133 (w1444) @(2371, 1500) /w:[ 46 45 76 -1 ]
  HD g263 (.B(w1254), .A(A1), .CrIn(w1347), .PrIn(w1444), .PrOut(w1349), .BOut(w1350), .Q(w1351), .CrOut(Cr29));   //: @(3342, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>65 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g68 (.B(w84), .A(w81), .CrIn(w312), .PrIn(w307), .PrOut(w313), .BOut(w314), .Q(w470), .CrOut(w306));   //: @(937, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  //: IN g31 (A) @(1274,-297) /sn:0 /R:2 /w:[ 0 ]
  HD g22 (.B(w42), .A(w62), .CrIn(w72), .PrIn(w73), .PrOut(w74), .BOut(w296), .Q(w346), .CrOut(w77));   //: @(-503, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g225 (.B(w1051), .A(w1011), .CrIn(w1130), .PrIn(w1105), .PrOut(w1126), .BOut(w1147), .Q(w1220), .CrOut(Cr26));   //: @(585, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g283 (.B(w1456), .A(w1351), .CrIn(w1458), .PrIn(w1445), .PrOut(w1459), .BOut(w1460), .Q(w1461), .CrOut(w1443));   //: @(3342, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  NandNOT g87 (.in1(w412), .out(w413));   //: @(-1340, 851) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  NandNOT g231 (.in1(w1180), .out(w1181));   //: @(159, 2090) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  assign A4 = A[4]; //: TAP g317 @(1163,-299) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  HD g83 (.B(w294), .A(A11), .CrIn(w387), .PrIn(w1444), .PrOut(w389), .BOut(w390), .Q(w391), .CrOut(w0));   //: @(1470, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>85 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g328 (w1444) @(-283, 129) /w:[ 18 -1 17 104 ]
  HD g41 (.B(B13), .A(w1444), .CrIn(w146), .PrIn(w141), .PrOut(w147), .BOut(w148), .Q(w149), .CrOut(w140));   //: @(-1604, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>119 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g203 (.B(w942), .A(w948), .CrIn(w989), .PrIn(w1037), .PrOut(w988), .BOut(w1131), .Q(w1039), .CrOut(w1040));   //: @(-134, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g264 (.B(w1261), .A(w1304), .CrIn(w1354), .PrIn(w1355), .PrOut(w1356), .BOut(w1493), .Q(w1498), .CrOut(w1359));   //: @(1664, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g42 (.B(B14), .A(w1444), .CrIn(w137), .PrIn(w147), .PrOut(w133), .BOut(w153), .Q(w154), .CrOut(w146));   //: @(-1786, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g138 (.B(w680), .A(w681), .CrIn(w682), .PrIn(w683), .PrOut(w684), .BOut(w685), .Q(w686), .CrOut(w687));   //: @(418, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  NandNOT g213 (.in1(w1084), .out(w1085));   //: @(-29, 1937) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: joint g151 (w1444) @(2564, 1647) /w:[ 48 47 74 -1 ]
  HD g293 (.B(w1515), .A(w1428), .CrIn(w1469), .PrIn(w1517), .PrOut(w1468), .BOut(w1518), .Q(w1519), .CrOut(w1520));   //: @(758, 2518) /sz:(123, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g66 (.B(w296), .A(w297), .CrIn(w298), .PrIn(w299), .PrOut(w300), .BOut(w392), .Q(w442), .CrOut(w303));   //: @(-318, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g167 (.B(w843), .A(w756), .CrIn(w797), .PrIn(w845), .PrOut(w796), .BOut(w846), .Q(w847), .CrOut(w848));   //: @(-503, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g146 (.B(w635), .A(w590), .CrIn(w724), .PrIn(w684), .PrOut(w720), .BOut(w825), .Q(w732), .CrOut(w682));   //: @(234, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g153 (.B(w667), .A(w762), .CrIn(w746), .PrIn(w721), .PrOut(w742), .BOut(w763), .Q(w836), .CrOut(Cr18));   //: @(-134, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g162 (.B(w814), .A(w732), .CrIn(Cr20), .PrIn(w816), .PrOut(w817), .BOut(w910), .Q(w954), .CrOut(w820));   //: @(234, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  //: joint g241 (w1444) @(3496, 2404) /w:[ 58 57 64 -1 ]
  assign A3 = A[3]; //: TAP g318 @(1186,-299) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign A13 = A[13]; //: TAP g34 @(990,-299) /sn:0 /R:1 /w:[ 1 28 27 ] /ss:1
  HD g46 (.B(w148), .A(w143), .CrIn(w185), .PrIn(w186), .PrOut(w187), .BOut(w188), .Q(w189), .CrOut(w190));   //: @(-1420, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  //: joint g5 (w1444) @(1099, 363) /w:[ 32 31 90 -1 ]
  HD g118 (.B(w573), .A(w574), .CrIn(w517), .PrIn(w544), .PrOut(w513), .BOut(w669), .Q(w576), .CrOut(w543));   //: @(585, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g84 (.B(w392), .A(w344), .CrIn(w394), .PrIn(w395), .PrOut(w396), .BOut(w397), .Q(w538), .CrOut(w399));   //: @(-134, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g112 (.B(w456), .A(w548), .CrIn(w549), .PrIn(w550), .PrOut(w551), .BOut(w552), .Q(w658), .CrOut(w554));   //: @(-688, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g201 (.B(w1021), .A(w908), .CrIn(w1023), .PrIn(w1002), .PrOut(w1024), .BOut(w1117), .Q(w1150), .CrOut(w1000));   //: @(1664, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  //: joint g61 (w1444) @(1634, 861) /w:[ 38 37 84 -1 ]
  HD g279 (.B(w1339), .A(w1434), .CrIn(w1418), .PrIn(w1393), .PrOut(w1414), .BOut(w1529), .Q(w1508), .CrOut(Cr32));   //: @(1108, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g21 (.B(w37), .A(A13), .CrIn(w67), .PrIn(w1444), .PrOut(w69), .BOut(w70), .Q(w71), .CrOut(Cr5));   //: @(1108, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>89 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g255 (.B(w1309), .A(w1310), .CrIn(w1311), .PrIn(w1290), .PrOut(w1312), .BOut(w1313), .Q(w1438), .CrOut(w1288));   //: @(2211, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  assign A15 = A[15]; //: TAP g32 @(955,-299) /sn:0 /R:1 /w:[ 1 32 31 ] /ss:1
  assign B4 = B[4]; //: TAP g295 @(753,-300) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  HD g20 (.B(w1), .A(w16), .CrIn(w55), .PrIn(w50), .PrOut(w54), .BOut(w65), .Q(w66), .CrOut(w49));   //: @(418, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g97 (w1444) @(1278, 529) /w:[ 34 33 88 -1 ]
  assign A10 = A[10]; //: TAP g311 @(1047,-299) /sn:0 /R:1 /w:[ 1 22 21 ] /ss:1
  HD g134 (.B(w661), .A(w507), .CrIn(w621), .PrIn(w601), .PrOut(w617), .BOut(w663), .Q(w664), .CrOut(w600));   //: @(1290, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g175 (.B(w788), .A(w775), .CrIn(w882), .PrIn(w869), .PrOut(w883), .BOut(w884), .Q(w885), .CrOut(w867));   //: @(2211, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g176 (.B(w794), .A(w789), .CrIn(w888), .PrIn(w883), .PrOut(w889), .BOut(w982), .Q(w891), .CrOut(w882));   //: @(2034, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g240 (.B(w1139), .A(w1129), .CrIn(w1232), .PrIn(w1223), .PrOut(w1229), .BOut(w1235), .Q(w1236), .CrOut(w1221));   //: @(418, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g89 (.B(w422), .A(w423), .CrIn(w424), .PrIn(w425), .PrOut(w426), .BOut(w427), .Q(w428), .CrOut(w429));   //: @(761, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  NandNOT g15 (.in1(w53), .out(w156));   //: @(-1885, 350) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g148 (.B(w648), .A(w740), .CrIn(w741), .PrIn(w742), .PrOut(w743), .BOut(w744), .Q(w745), .CrOut(w746));   //: @(-318, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g147 (.B(w733), .A(w620), .CrIn(w735), .PrIn(w714), .PrOut(w736), .BOut(w829), .Q(w862), .CrOut(w712));   //: @(1108, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g165 (.B(w829), .A(w716), .CrIn(w831), .PrIn(w810), .PrOut(w832), .BOut(w925), .Q(w834), .CrOut(w808));   //: @(1290, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g247 (.B(w1172), .A(w1265), .CrIn(w1266), .PrIn(w1253), .PrOut(w1267), .BOut(w1268), .Q(w1367), .CrOut(w1251));   //: @(2965, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g252 (.B(w1202), .A(w1212), .CrIn(Cr30), .PrIn(w1296), .PrOut(w1297), .BOut(w1390), .Q(w1434), .CrOut(w1300));   //: @(1108, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g336 (w1444) @(-1751, 129) /w:[ 2 -1 120 1 ]
  HD g62 (.B(w65), .A(w52), .CrIn(w237), .PrIn(w83), .PrOut(w233), .BOut(w279), .Q(w327), .CrOut(w82));   //: @(585, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g160 (.B(w707), .A(w799), .CrIn(w800), .PrIn(w801), .PrOut(w802), .BOut(w803), .Q(w918), .CrOut(w805));   //: @(937, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g218 (.B(w1019), .A(w974), .CrIn(w1108), .PrIn(w1068), .PrOut(w1104), .BOut(w1115), .Q(w1199), .CrOut(w1066));   //: @(937, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g55 (.B(w61), .A(w163), .CrIn(w77), .PrIn(w226), .PrOut(w73), .BOut(w247), .Q(w297), .CrOut(w224));   //: @(-318, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  NandNOT g195 (.in1(w988), .out(w989));   //: @(-213, 1788) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g53 (.B(w169), .A(w66), .CrIn(w232), .PrIn(w233), .PrOut(w234), .BOut(w326), .Q(w350), .CrOut(w237));   //: @(418, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g13 (.B(w17), .A(w24), .CrIn(w45), .PrIn(w34), .PrOut(w46), .BOut(w47), .Q(w218), .CrOut(w33));   //: @(761, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g135 (.B(w665), .A(w531), .CrIn(w650), .PrIn(w625), .PrOut(w646), .BOut(w667), .Q(w740), .CrOut(Cr16));   //: @(-318, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g139 (.B(w596), .A(w583), .CrIn(w690), .PrIn(w677), .PrOut(w691), .BOut(w784), .Q(w791), .CrOut(w675));   //: @(1858, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  assign B14 = B[14]; //: TAP g308 @(507,-300) /sn:0 /R:1 /w:[ 1 30 29 ] /ss:1
  HD g116 (.B(w471), .A(w566), .CrIn(w525), .PrIn(w505), .PrOut(w521), .BOut(w661), .Q(w615), .CrOut(w504));   //: @(1108, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g4 (.B(B0), .A(A15), .CrIn(w23), .PrIn(w1444), .PrOut(w19), .BOut(w28), .Q(w24), .CrOut(Cr3));   //: @(761, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>93 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g246 (.B(w1165), .A(w1257), .CrIn(w1258), .PrIn(w1259), .PrOut(w1260), .BOut(w1261), .Q(w1262), .CrOut(w1263));   //: @(1470, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g157 (.B(w784), .A(w785), .CrIn(w786), .PrIn(w773), .PrOut(w787), .BOut(w788), .Q(w789), .CrOut(w771));   //: @(2034, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g197 (.B(w998), .A(w952), .CrIn(w1000), .PrIn(w1001), .PrOut(w1002), .BOut(w1094), .Q(w1004), .CrOut(w1005));   //: @(1858, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g271 (.B(w1397), .A(w1284), .CrIn(w1359), .PrIn(w1378), .PrOut(w1355), .BOut(w1399), .Q(w1449), .CrOut(w1376));   //: @(1858, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g17 (.B(w29), .A(w129), .CrIn(w44), .PrIn(w161), .PrOut(w40), .BOut(w61), .Q(w62), .CrOut(w159));   //: @(-503, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g137 (.B(w582), .A(A8), .CrIn(w675), .PrIn(w1444), .PrOut(w677), .BOut(w769), .Q(w785), .CrOut(Cr17));   //: @(2034, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>79 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g280 (.B(w1437), .A(w1438), .CrIn(w1381), .PrIn(w1408), .PrOut(w1377), .BOut(w1439), .Q(w1471), .CrOut(w1407));   //: @(2211, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  //: joint g326 (w1444) @(89, 129) /w:[ 22 -1 21 100 ]
  HD g282 (.B(w1493), .A(w1449), .CrIn(w1450), .PrIn(w1451), .PrOut(w1452), .BOut(w1453), .Q(w1454), .CrOut(w1455));   //: @(1858, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g77 (.B(w270), .A(w364), .CrIn(w317), .PrIn(w365), .PrOut(w316), .BOut(w459), .Q(w367), .CrOut(w368));   //: @(-1420, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g214 (.B(w995), .A(w1056), .CrIn(w1088), .PrIn(w1089), .PrOut(w1090), .BOut(w1182), .Q(w1092), .CrOut(w1093));   //: @(1470, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g327 (w1444) @(-99, 129) /w:[ 20 -1 19 102 ]
  HD g291 (.B(w1409), .A(w1502), .CrIn(w1503), .PrIn(w1482), .PrOut(w1504), .BOut(w1505), .Q(w1506), .CrOut(w1480));   //: @(2592, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g275 (.B(w1419), .A(w1420), .CrIn(w1373), .PrIn(w1421), .PrOut(w1372), .BOut(w1515), .Q(w1423), .CrOut(w1424));   //: @(588, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  NandNOT g51 (.in1(w220), .out(w221));   //: @(-1701, 516) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g144 (.B(w718), .A(w719), .CrIn(Cr18), .PrIn(w720), .PrOut(w721), .BOut(w814), .Q(w723), .CrOut(w724));   //: @(54, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g259 (w1444) @(3667, 2550) /w:[ 60 59 62 -1 ]
  HD g161 (.B(w806), .A(w760), .CrIn(w808), .PrIn(w809), .PrOut(w810), .BOut(w811), .Q(w926), .CrOut(w813));   //: @(1470, 1468) /sz:(122, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g190 (.B(w863), .A(w834), .CrIn(w901), .PrIn(w928), .PrOut(w897), .BOut(w1053), .Q(w991), .CrOut(w927));   //: @(1290, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g296 (.B(w1525), .A(w1526), .CrIn(w1485), .PrIn(w1465), .PrOut(w1481), .BOut(w1527), .Q(w1528), .CrOut(w1464));   //: @(2965, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g103 (.B(w496), .A(w391), .CrIn(w498), .PrIn(w485), .PrOut(w499), .BOut(w500), .Q(w501), .CrOut(w483));   //: @(1470, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g65 (.B(w70), .A(A12), .CrIn(w291), .PrIn(w1444), .PrOut(w293), .BOut(w294), .Q(w308), .CrOut(Cr9));   //: @(1290, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>87 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  assign B10 = B[10]; //: TAP g304 @(615,-300) /sn:0 /R:1 /w:[ 1 22 21 ] /ss:1
  HD g72 (.B(w242), .A(w335), .CrIn(Cr10), .PrIn(w336), .PrOut(w337), .BOut(w338), .Q(w339), .CrOut(w340));   //: @(-688, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g185 (.B(w846), .A(w852), .CrIn(w893), .PrIn(w941), .PrOut(w892), .BOut(w942), .Q(w943), .CrOut(w944));   //: @(-318, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g6 (w1444) @(2018, 1190) /w:[ 42 41 80 -1 ]
  HD g136 (.B(w669), .A(w670), .CrIn(w613), .PrIn(w640), .PrOut(w609), .BOut(w765), .Q(w703), .CrOut(w639));   //: @(761, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g142 (.B(w702), .A(w703), .CrIn(w704), .PrIn(w705), .PrOut(w706), .BOut(w707), .Q(w822), .CrOut(w709));   //: @(761, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g251 (.B(w1286), .A(w1287), .CrIn(w1288), .PrIn(w1289), .PrOut(w1290), .BOut(w1291), .Q(w1292), .CrOut(w1293));   //: @(2397, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: GROUND g277 (w1444) @(3705,2562) /sn:0 /w:[ 61 ]
  HD g124 (.B(w515), .A(w576), .CrIn(w608), .PrIn(w609), .PrOut(w610), .BOut(w702), .Q(w726), .CrOut(w613));   //: @(585, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g58 (.B(w188), .A(w206), .CrIn(w261), .PrIn(w262), .PrOut(w263), .BOut(w355), .Q(w370), .CrOut(w266));   //: @(-1238, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g56 (.B(w63), .A(w43), .CrIn(w244), .PrIn(w74), .PrOut(w240), .BOut(w345), .Q(w335), .CrOut(w72));   //: @(-688, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g7 (.B(B8), .A(w1444), .CrIn(w26), .PrIn(w127), .PrOut(w21), .BOut(w29), .Q(w27), .CrOut(w126));   //: @(-688, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>109 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g297 (.B(w1529), .A(w1530), .CrIn(w1514), .PrIn(w1489), .PrOut(w1510), .BOut(w1531), .Q(w1532), .CrOut(Cr34));   //: @(1290, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g98 (.B(w469), .A(w470), .CrIn(w429), .PrIn(w409), .PrOut(w425), .BOut(w471), .Q(w519), .CrOut(w408));   //: @(937, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g200 (.B(w1017), .A(w1018), .CrIn(w1012), .PrIn(w972), .PrOut(w1008), .BOut(w1019), .Q(w1020), .CrOut(w970));   //: @(761, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g229 (.B(w1076), .A(w1063), .CrIn(w1170), .PrIn(w1157), .PrOut(w1171), .BOut(w1172), .Q(w1173), .CrOut(w1155));   //: @(2781, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g204 (.B(w1041), .A(w1042), .CrIn(w1040), .PrIn(w1031), .PrOut(w1037), .BOut(w1043), .Q(w1132), .CrOut(w1029));   //: @(54, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g208 (.B(w1053), .A(w1054), .CrIn(w997), .PrIn(w1024), .PrOut(w993), .BOut(w1055), .Q(w1056), .CrOut(w1023));   //: @(1470, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g81 (.B(w377), .A(w378), .CrIn(w362), .PrIn(w337), .PrOut(w358), .BOut(w379), .Q(w452), .CrOut(Cr10));   //: @(-872, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g52 (.B(w162), .A(w223), .CrIn(w224), .PrIn(w225), .PrOut(w226), .BOut(w227), .Q(w228), .CrOut(w229));   //: @(-134, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g40 (.B(B15), .A(w1444), .CrIn(w104), .PrIn(w133), .PrOut(w4), .BOut(w135), .Q(w136), .CrOut(w137));   //: @(-1970, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>121 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  assign A8 = A[8]; //: TAP g313 @(1082,-299) /sn:0 /R:1 /w:[ 1 18 17 ] /ss:1
  //: joint g332 (w1444) @(-1021, 129) /w:[ 10 -1 9 112 ]
  HD g108 (.B(w526), .A(w527), .CrIn(Cr14), .PrIn(w528), .PrOut(w529), .BOut(w622), .Q(w531), .CrOut(w532));   //: @(-318, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g210 (.B(w1064), .A(w1065), .CrIn(w1066), .PrIn(w1067), .PrOut(w1068), .BOut(w1069), .Q(w1210), .CrOut(w1071));   //: @(1108, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  //: joint g330 (w1444) @(-653, 129) /w:[ 14 -1 13 108 ]
  HD g131 (.B(w651), .A(w652), .CrIn(w605), .PrIn(w653), .PrOut(w604), .BOut(w654), .Q(w655), .CrOut(w656));   //: @(-872, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  assign B5 = B[5]; //: TAP g299 @(733,-300) /sn:0 /R:1 /w:[ 1 12 11 ] /ss:1
  HD g290 (.B(w1497), .A(w1498), .CrIn(w1492), .PrIn(w1452), .PrOut(w1488), .BOut(w1499), .Q(w1500), .CrOut(w1450));   //: @(1664, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g266 (.B(w1274), .A(w1367), .CrIn(w1368), .PrIn(w1363), .PrOut(w1369), .BOut(w1370), .Q(w1526), .CrOut(w1362));   //: @(2965, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g96 (.B(w465), .A(w466), .CrIn(w464), .PrIn(w455), .PrOut(w461), .BOut(w561), .Q(w468), .CrOut(w453));   //: @(-1056, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g209 (.B(w1057), .A(A4), .CrIn(w1059), .PrIn(w1444), .PrOut(w1061), .BOut(w1062), .Q(w1063), .CrOut(Cr23));   //: @(2781, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>71 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g294 (.B(w1521), .A(w1417), .CrIn(w1520), .PrIn(w1511), .PrOut(w1517), .BOut(w1523), .Q(w1524), .CrOut(w1509));   //: @(937, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g117 (.B(w569), .A(w570), .CrIn(w554), .PrIn(w529), .PrOut(w550), .BOut(w665), .Q(w644), .CrOut(Cr14));   //: @(-503, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g221 (.B(w1131), .A(w1132), .CrIn(w1085), .PrIn(w1133), .PrOut(w1084), .BOut(w1134), .Q(w1135), .CrOut(w1136));   //: @(54, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  assign A6 = A[6]; //: TAP g315 @(1121,-299) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  HD g78 (.B(w369), .A(w370), .CrIn(w368), .PrIn(w359), .PrOut(w365), .BOut(w465), .Q(w372), .CrOut(w357));   //: @(-1238, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g223 (w1444) @(3310, 2250) /w:[ 56 55 66 -1 ]
  HD g113 (.B(w555), .A(w468), .CrIn(w509), .PrIn(w557), .PrOut(w508), .BOut(w651), .Q(w559), .CrOut(w560));   //: @(-1056, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  NandNOT g105 (.in1(w508), .out(w509));   //: @(-1149, 1019) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g155 (.B(w769), .A(A7), .CrIn(w771), .PrIn(w1444), .PrOut(w773), .BOut(w774), .Q(w775), .CrOut(w80));   //: @(2211, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>77 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g219 (.B(w1117), .A(w1004), .CrIn(w1119), .PrIn(w1098), .PrOut(w1120), .BOut(w1213), .Q(w1122), .CrOut(w1096));   //: @(1858, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  //: joint g205 (w1444) @(3122, 2102) /w:[ 54 53 68 -1 ]
  assign B9 = B[9]; //: TAP g303 @(640,-300) /sn:0 /R:1 /w:[ 1 20 19 ] /ss:1
  HD g292 (.B(w1507), .A(w1508), .CrIn(w1509), .PrIn(w1510), .PrOut(w1511), .BOut(w1512), .Q(w1513), .CrOut(w1514));   //: @(1108, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g43 (.B(w128), .A(w123), .CrIn(w159), .PrIn(w160), .PrOut(w161), .BOut(w162), .Q(w163), .CrOut(w164));   //: @(-318, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g38 (.B(B12), .A(w1444), .CrIn(w140), .PrIn(w14), .PrOut(w141), .BOut(w142), .Q(w143), .CrOut(Cr6));   //: @(-1420, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>117 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g212 (.B(w986), .A(w1079), .CrIn(w1080), .PrIn(w1075), .PrOut(w1081), .BOut(w1174), .Q(w1238), .CrOut(w1074));   //: @(2397, 1919) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  assign A0 = A[0]; //: TAP g321 @(1258,-299) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  assign B11 = B[11]; //: TAP g305 @(588,-300) /sn:0 /R:1 /w:[ 1 24 23 ] /ss:1
  HD g287 (.B(w1387), .A(w1479), .CrIn(w1480), .PrIn(w1481), .PrOut(w1482), .BOut(w1483), .Q(w1484), .CrOut(w1485));   //: @(2781, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g48 (.B(w153), .A(w149), .CrIn(w196), .PrIn(w187), .PrOut(w193), .BOut(w199), .Q(w200), .CrOut(w185));   //: @(-1604, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  assign A2 = A[2]; //: TAP g319 @(1212,-299) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  HD g276 (.B(w1331), .A(w1426), .CrIn(w1424), .PrIn(w1415), .PrOut(w1421), .BOut(w1521), .Q(w1428), .CrOut(w1413));   //: @(761, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g237 (.B(w1213), .A(w1100), .CrIn(w1215), .PrIn(w1194), .PrOut(w1216), .BOut(w1309), .Q(w1342), .CrOut(w1192));   //: @(2034, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g122 (.B(w506), .A(w501), .CrIn(w600), .PrIn(w595), .PrOut(w601), .BOut(w602), .Q(w603), .CrOut(w594));   //: @(1470, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  //: joint g322 (w1444) @(928, 190) /w:[ 30 29 92 -1 ]
  HD g80 (.B(w279), .A(w374), .CrIn(w333), .PrIn(w313), .PrOut(w329), .BOut(w469), .Q(w423), .CrOut(w312));   //: @(761, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g95 (.B(w459), .A(w372), .CrIn(w413), .PrIn(w461), .PrOut(w412), .BOut(w555), .Q(w463), .CrOut(w464));   //: @(-1238, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g170 (.B(w853), .A(w699), .CrIn(w813), .PrIn(w793), .PrOut(w809), .BOut(w949), .Q(w856), .CrOut(w792));   //: @(1664, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g178 (.B(w803), .A(w864), .CrIn(w896), .PrIn(w897), .PrOut(w898), .BOut(w899), .Q(w1014), .CrOut(w901));   //: @(1108, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g189 (.B(w859), .A(w954), .CrIn(w938), .PrIn(w913), .PrOut(w934), .BOut(w1049), .Q(w956), .CrOut(Cr22));   //: @(234, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g324 (w1444) @(453, 129) /w:[ 26 -1 25 96 ]
  HD g269 (.B(w1291), .A(w1383), .CrIn(w1384), .PrIn(w1385), .PrOut(w1386), .BOut(w1387), .Q(w1502), .CrOut(w1389));   //: @(2592, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g182 (.B(w827), .A(w922), .CrIn(w916), .PrIn(w876), .PrOut(w912), .BOut(w1017), .Q(w924), .CrOut(w874));   //: @(585, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g335 (w1444) @(-1569, 129) /w:[ 4 -1 3 118 ]
  HD g90 (.B(w338), .A(w348), .CrIn(Cr12), .PrIn(w432), .PrOut(w433), .BOut(w526), .Q(w570), .CrOut(w436));   //: @(-503, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g268 (.B(w1374), .A(w1375), .CrIn(w1376), .PrIn(w1377), .PrOut(w1378), .BOut(w1470), .Q(w1380), .CrOut(w1381));   //: @(2034, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g128 (.B(w539), .A(w634), .CrIn(w628), .PrIn(w588), .PrOut(w624), .BOut(w635), .Q(w719), .CrOut(w586));   //: @(54, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g2 (.B(B2), .A(w1444), .CrIn(w7), .PrIn(w11), .PrOut(w3), .BOut(w8), .Q(w16), .CrOut(w15));   //: @(418, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>97 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g174 (.B(w872), .A(w873), .CrIn(w874), .PrIn(w875), .PrOut(w876), .BOut(w968), .Q(w1018), .CrOut(w879));   //: @(761, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g91 (.B(w343), .A(w438), .CrIn(w399), .PrIn(w418), .PrOut(w395), .BOut(w533), .Q(w489), .CrOut(w416));   //: @(54, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  NandNOT g285 (.in1(w1468), .out(w1469));   //: @(660, 2532) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g265 (.B(w1268), .A(w1361), .CrIn(w1362), .PrIn(w1349), .PrOut(w1363), .BOut(w1456), .Q(w1365), .CrOut(w1347));   //: @(3149, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  NandNOT g141 (.in1(w700), .out(w701));   //: @(-772, 1337) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: OUT g338 (Q) @(4164,2507) /sn:0 /w:[ 0 ]
  assign B2 = B[2]; //: TAP g29 @(797,-300) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  HD g288 (.B(w1486), .A(w1404), .CrIn(Cr34), .PrIn(w1488), .PrOut(w1489), .BOut(w1490), .Q(w1491), .CrOut(w1492));   //: @(1470, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g278 (.B(w1335), .A(w1430), .CrIn(w1389), .PrIn(w1369), .PrOut(w1385), .BOut(w1525), .Q(w1479), .CrOut(w1368));   //: @(2781, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g168 (.B(w755), .A(w745), .CrIn(w848), .PrIn(w839), .PrOut(w845), .BOut(w851), .Q(w852), .CrOut(w837));   //: @(-318, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<0 Ro0<0 ]
  HD g18 (.B(w13), .A(w31), .CrIn(w60), .PrIn(w41), .PrOut(w56), .BOut(w63), .Q(w64), .CrOut(w39));   //: @(-872, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g199 (.B(w919), .A(w1014), .CrIn(w975), .PrIn(w994), .PrOut(w971), .BOut(w1109), .Q(w1065), .CrOut(w992));   //: @(1108, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g119 (.B(w577), .A(A9), .CrIn(w579), .PrIn(w1444), .PrOut(w581), .BOut(w582), .Q(w583), .CrOut(w20));   //: @(1858, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>81 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g329 (w1444) @(-468, 129) /w:[ 16 -1 15 106 ]
  HD g154 (.B(w765), .A(w766), .CrIn(w709), .PrIn(w736), .PrOut(w705), .BOut(w861), .Q(w799), .CrOut(w735));   //: @(937, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g173 (.B(w774), .A(A6), .CrIn(w867), .PrIn(w1444), .PrOut(w869), .BOut(w961), .Q(w871), .CrOut(Cr21));   //: @(2397, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>75 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g172 (.B(w861), .A(w862), .CrIn(w805), .PrIn(w832), .PrOut(w801), .BOut(w863), .Q(w864), .CrOut(w831));   //: @(1108, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  HD g184 (.B(w840), .A(w932), .CrIn(w933), .PrIn(w934), .PrOut(w935), .BOut(w1027), .Q(w1042), .CrOut(w938));   //: @(54, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  HD g188 (.B(w949), .A(w795), .CrIn(w909), .PrIn(w889), .PrOut(w905), .BOut(w1045), .Q(w952), .CrOut(w888));   //: @(1858, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g256 (.B(w1315), .A(w1244), .CrIn(w1317), .PrIn(w1318), .PrOut(w1319), .BOut(w1320), .Q(w1426), .CrOut(w1322));   //: @(761, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g261 (.B(w1243), .A(w1338), .CrIn(w1322), .PrIn(w1297), .PrOut(w1318), .BOut(w1339), .Q(w1412), .CrOut(Cr30));   //: @(937, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g50 (.B(w122), .A(w117), .CrIn(w164), .PrIn(w180), .PrOut(w160), .BOut(w285), .Q(w223), .CrOut(w179));   //: @(-134, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  HD g193 (.B(w884), .A(w871), .CrIn(w978), .PrIn(w965), .PrOut(w979), .BOut(w1072), .Q(w1079), .CrOut(w963));   //: @(2397, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g73 (.B(w247), .A(w228), .CrIn(w303), .PrIn(w322), .PrOut(w299), .BOut(w343), .Q(w344), .CrOut(w320));   //: @(-134, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g9 (.B(B10), .A(w1444), .CrIn(w10), .PrIn(w12), .PrOut(w6), .BOut(w13), .Q(w32), .CrOut(w22));   //: @(-1056, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>113 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  //: joint g169 (w1444) @(2763, 1800) /w:[ 50 49 72 -1 ]
  HD g102 (.B(w397), .A(w489), .CrIn(w490), .PrIn(w491), .PrOut(w492), .BOut(w584), .Q(w634), .CrOut(w495));   //: @(54, 999) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g71 (.B(w326), .A(w327), .CrIn(w328), .PrIn(w329), .PrOut(w330), .BOut(w422), .Q(w332), .CrOut(w333));   //: @(585, 660) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g59 (.B(w194), .A(w200), .CrIn(w221), .PrIn(w269), .PrOut(w220), .BOut(w270), .Q(w271), .CrOut(w272));   //: @(-1604, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g186 (.B(w851), .A(w841), .CrIn(w944), .PrIn(w935), .PrOut(w941), .BOut(w1041), .Q(w948), .CrOut(w933));   //: @(-134, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  NandNOT g249 (.in1(w1276), .out(w1277));   //: @(345, 2236) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g99 (.B(w379), .A(w339), .CrIn(w458), .PrIn(w433), .PrOut(w454), .BOut(w569), .Q(w548), .CrOut(Cr12));   //: @(-688, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g180 (.B(w910), .A(w911), .CrIn(Cr22), .PrIn(w912), .PrOut(w913), .BOut(w1006), .Q(w915), .CrOut(w916));   //: @(418, 1615) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g45 (.B(w116), .A(w111), .CrIn(w179), .PrIn(w168), .PrOut(w180), .BOut(w253), .Q(w286), .CrOut(w167));   //: @(54, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g36 (.B(B5), .A(w1444), .CrIn(w114), .PrIn(w109), .PrOut(w115), .BOut(w116), .Q(w117), .CrOut(w107));   //: @(-134, 158) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>103 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<1 Ro0<1 ]
  NandNOT g69 (.in1(w316), .out(w317));   //: @(-1511, 679) /sz:(47, 62) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  HD g156 (.B(w685), .A(w777), .CrIn(w778), .PrIn(w779), .PrOut(w780), .BOut(w872), .Q(w922), .CrOut(w783));   //: @(585, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g254 (.B(w1211), .A(w1166), .CrIn(w1300), .PrIn(w1260), .PrOut(w1296), .BOut(w1307), .Q(w1391), .CrOut(w1258));   //: @(1290, 2218) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  assign Q = {Cr3, Cr4, Cr5, Cr9, w0, Cr13, w20, Cr17, w80, Cr21, w86, Cr23, Cr27, w89, Cr29, Cr31}; //: CONCAT g337  @(4100,2507) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: joint g325 (w1444) @(269, 129) /w:[ 24 -1 23 98 ]
  assign A1 = A[1]; //: TAP g320 @(1237,-299) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  HD g273 (.B(w1313), .A(w1292), .CrIn(w1407), .PrIn(w1386), .PrOut(w1408), .BOut(w1409), .Q(w1410), .CrOut(w1384));   //: @(2397, 2372) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g191 (.B(w961), .A(A5), .CrIn(w963), .PrIn(w1444), .PrOut(w965), .BOut(w1057), .Q(w1073), .CrOut(w86));   //: @(2592, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>73 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g232 (.B(w1182), .A(w1152), .CrIn(w1184), .PrIn(w1185), .PrOut(w1186), .BOut(w1278), .Q(w1302), .CrOut(w1189));   //: @(1664, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g233 (.B(w1190), .A(w1191), .CrIn(w1192), .PrIn(w1193), .PrOut(w1194), .BOut(w1286), .Q(w1310), .CrOut(w1197));   //: @(2211, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  assign B1 = B[1]; //: TAP g28 @(819,-300) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  HD g286 (.B(w1470), .A(w1471), .CrIn(w1472), .PrIn(w1473), .PrOut(w1474), .BOut(w1475), .Q(w1476), .CrOut(w1477));   //: @(2211, 2518) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g57 (.B(w253), .A(w170), .CrIn(w255), .PrIn(w234), .PrOut(w256), .BOut(w349), .Q(w382), .CrOut(w232));   //: @(234, 497) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>0 Lo0<0 Bo0<0 Bo1<0 Ro0<1 ]
  HD g239 (.B(w1134), .A(w1228), .CrIn(w1181), .PrIn(w1229), .PrOut(w1180), .BOut(w1323), .Q(w1231), .CrOut(w1232));   //: @(234, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g242 (.B(w1237), .A(w1238), .CrIn(w1197), .PrIn(w1177), .PrOut(w1193), .BOut(w1239), .Q(w1287), .CrOut(w1176));   //: @(2397, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g14 (.B(w8), .A(w25), .CrIn(w49), .PrIn(w46), .PrOut(w50), .BOut(w217), .Q(w52), .CrOut(w45));   //: @(585, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g11 (.B(w28), .A(A14), .CrIn(w33), .PrIn(w1444), .PrOut(w34), .BOut(w37), .Q(w38), .CrOut(Cr4));   //: @(937, 331) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>91 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g150 (.B(w659), .A(w649), .CrIn(w752), .PrIn(w743), .PrOut(w749), .BOut(w755), .Q(w756), .CrOut(w741));   //: @(-503, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Ro0<0 ]
  //: joint g333 (w1444) @(-1203, 129) /w:[ 8 -1 7 114 ]
  //: joint g187 (w1444) @(2955, 1951) /w:[ 52 51 70 -1 ]
  NandNOT g123 (.in1(w604), .out(w605));   //: @(-951, 1176) /sz:(47, 63) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  //: joint g79 (w1444) @(1453, 692) /w:[ 36 35 86 -1 ]
  //: joint g115 (w1444) @(2204, 1348) /w:[ 44 43 78 -1 ]
  HD g145 (.B(w631), .A(w726), .CrIn(w687), .PrIn(w706), .PrOut(w683), .BOut(w821), .Q(w777), .CrOut(w704));   //: @(585, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<0 Bo1<0 Ro0<0 ]
  HD g235 (.B(w1111), .A(w1092), .CrIn(w1167), .PrIn(w1186), .PrOut(w1163), .BOut(w1207), .Q(w1257), .CrOut(w1184));   //: @(1470, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]
  HD g129 (.B(w545), .A(w638), .CrIn(w639), .PrIn(w618), .PrOut(w640), .BOut(w733), .Q(w766), .CrOut(w616));   //: @(937, 1158) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<0 Ro0<1 ]
  HD g236 (.B(w1115), .A(w1210), .CrIn(w1204), .PrIn(w1164), .PrOut(w1200), .BOut(w1211), .Q(w1212), .CrOut(w1162));   //: @(1108, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Ro0<0 ]
  assign B0 = B[0]; //: TAP g27 @(837,-300) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  HD g202 (.B(w1027), .A(w956), .CrIn(w1029), .PrIn(w1030), .PrOut(w1031), .BOut(w1032), .Q(w1033), .CrOut(w1034));   //: @(234, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  HD g227 (.B(w1062), .A(A3), .CrIn(w1155), .PrIn(w1444), .PrOut(w1157), .BOut(w1158), .Q(w1265), .CrOut(Cr27));   //: @(2965, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>69 Lo0<1 Bo0<0 Bo1<1 Ro0<0 ]
  HD g171 (.B(w763), .A(w723), .CrIn(w842), .PrIn(w817), .PrOut(w838), .BOut(w859), .Q(w932), .CrOut(Cr20));   //: @(54, 1468) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g88 (.B(w323), .A(w415), .CrIn(w416), .PrIn(w417), .PrOut(w418), .BOut(w419), .Q(w534), .CrOut(w421));   //: @(234, 829) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Ro0<0 ]
  HD g238 (.B(w1128), .A(w1220), .CrIn(w1221), .PrIn(w1222), .PrOut(w1223), .BOut(w1315), .Q(w1225), .CrOut(w1226));   //: @(585, 2070) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>1 Ri0>0 Lo0<0 Bo0<1 Bo1<1 Ro0<1 ]
  assign A7 = A[7]; //: TAP g314 @(1101,-299) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  HD g140 (.B(w602), .A(w597), .CrIn(w696), .PrIn(w691), .PrOut(w697), .BOut(w790), .Q(w699), .CrOut(w690));   //: @(1664, 1316) /sz:(120, 103) /sn:0 /p:[ Ti0>0 Ti1>1 Li0>1 Ri0>1 Lo0<0 Bo0<0 Bo1<1 Ro0<0 ]
  HD g207 (.B(w1049), .A(w915), .CrIn(w1034), .PrIn(w1009), .PrOut(w1030), .BOut(w1051), .Q(w1052), .CrOut(Cr24));   //: @(418, 1768) /sz:(120, 103) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin HD
module HD(PrOut, PrIn, B, A, CrIn, Q, CrOut, BOut);
//: interface  /sz:(120, 103) /bd:[ Ti0>B(76/120) Ti1>A(35/120) Li0>CrIn(67/103) Ri0>PrIn(32/103) Lo0<PrOut(33/103) Bo0<BOut(84/120) Bo1<Q(37/120) Ro0<CrOut(64/103) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(294,151)(294,110){1}
//: {2}(296,108)(427,108)(427,134){3}
//: {4}(429,136)(444,136)(444,150){5}
//: {6}(425,136)(414,136)(414,150){7}
//: {8}(294,106)(294,86){9}
input PrIn;    //: /sn:0 {0}(361,135)(361,179)(333,179){1}
output Q;    //: /sn:0 {0}(232,319)(232,440)(233,440)(233,443){1}
input A;    //: /sn:0 {0}(199,269)(199,112)(253,112){1}
//: {2}(255,110)(255,87){3}
//: {4}(255,114)(255,151){5}
output PrOut;    //: /sn:0 {0}(89,182)(221,182){1}
output BOut;    //: /sn:0 {0}(426,443)(426,334)(426,334)(426,223){1}
input CrIn;    //: /sn:0 {0}(97,294)(119,294){1}
//: {2}(123,294)(168,294){3}
//: {4}(121,296)(121,309){5}
//: {6}(123,311)(135,311)(135,339){7}
//: {8}(119,311)(105,311)(105,339){9}
output CrOut;    //: /sn:0 {0}(122,443)(122,401){1}
wire w4;    //: /sn:0 {0}(272,269)(272,215){1}
//: enddecls

  //: joint g8 (A) @(255, 112) /w:[ -1 2 1 4 ]
  MUX g4 (.B(w4), .A(A), .Cin(CrIn), .Y(Q));   //: @(169, 270) /sz:(121, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Bo0<0 ]
  //: OUT g16 (PrOut) @(92,182) /sn:0 /R:2 /w:[ 0 ]
  //: IN g3 (PrIn) @(361,133) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (B) @(294,84) /sn:0 /R:3 /w:[ 9 ]
  //: IN g1 (A) @(255,85) /sn:0 /R:3 /w:[ 3 ]
  //: IN g10 (CrIn) @(95,294) /sn:0 /w:[ 0 ]
  //: joint g6 (B) @(294, 108) /w:[ 2 8 -1 1 ]
  //: OUT g9 (Q) @(233,440) /sn:0 /R:3 /w:[ 1 ]
  //: joint g7 (B) @(427, 136) /w:[ 4 3 6 -1 ]
  //: joint g12 (CrIn) @(121, 294) /w:[ 2 -1 1 4 ]
  //: joint g14 (CrIn) @(121, 311) /w:[ 6 5 8 -1 ]
  NandAND g11 (.in1(CrIn), .in2(CrIn), .out(CrOut));   //: @(85, 340) /sz:(64, 60) /R:3 /sn:0 /p:[ Ti0>7 Ti1>9 Bo0<1 ]
  NandAND g5 (.in1(B), .in2(B), .out(BOut));   //: @(400, 151) /sz:(58, 71) /R:3 /sn:0 /p:[ Ti0>7 Ti1>5 Bo0<1 ]
  //: OUT g15 (CrOut) @(122,440) /sn:0 /R:3 /w:[ 0 ]
  FS g0 (.A(A), .B(B), .PrIn(PrIn), .PrOut(PrOut), .D(w4));   //: @(222, 152) /sz:(110, 62) /sn:0 /p:[ Ti0>5 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  //: OUT g13 (BOut) @(426,440) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin RCA16
module RCA16(S, Cout, B, A);
//: interface  /sz:(89, 91) /bd:[ Ti0>A[15:0](23/89) Ti1>B[15:0](65/89) Lo0<Cout(41/91) Bo0<S[15:0](43/89) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [15:0] B;    //: /sn:0 {0}(#:1692,136)(1663,136){1}
//: {2}(1662,136)(1546,136){3}
//: {4}(1545,136)(1420,136){5}
//: {6}(1419,136)(1292,136){7}
//: {8}(1291,136)(1175,136){9}
//: {10}(1174,136)(1047,136){11}
//: {12}(1046,136)(923,136){13}
//: {14}(922,136)(806,136){15}
//: {16}(805,136)(688,136){17}
//: {18}(687,136)(556,136){19}
//: {20}(555,136)(425,136){21}
//: {22}(424,136)(309,136){23}
//: {24}(308,136)(181,136){25}
//: {26}(180,136)(55,136){27}
//: {28}(54,136)(-61,136){29}
//: {30}(-62,136)(-183,136){31}
//: {32}(-184,136)(-214,136){33}
input [15:0] A;    //: /sn:0 {0}(#:1650,189)(1627,189){1}
//: {2}(1626,189)(1506,189){3}
//: {4}(1505,189)(1380,189){5}
//: {6}(1379,189)(1252,189){7}
//: {8}(1251,189)(1135,189){9}
//: {10}(1134,189)(1007,189){11}
//: {12}(1006,189)(883,189){13}
//: {14}(882,189)(766,189){15}
//: {16}(765,189)(648,189){17}
//: {18}(647,189)(516,189){19}
//: {20}(515,189)(385,189){21}
//: {22}(384,189)(269,189){23}
//: {24}(268,189)(141,189){25}
//: {26}(140,189)(15,189){27}
//: {28}(14,189)(-101,189){29}
//: {30}(-102,189)(-223,189){31}
//: {32}(-224,189)(#:-250,189){33}
output Cout;    //: /sn:0 {0}(1794,512)(-293,512)(-293,281)(-244,281){1}
output [15:0] S;    //: /sn:0 {0}(#:1762,410)(1820,410){1}
wire w6;    //: /sn:0 {0}(269,193)(269,239){1}
wire w16;    //: /sn:0 {0}(141,193)(141,240){1}
wire w13;    //: /sn:0 {0}(-199,325)(-199,335)(1756,335){1}
wire w7;    //: /sn:0 {0}(364,276)(330,276){1}
wire w58;    //: /sn:0 {0}(709,273)(745,273){1}
wire w65;    //: /sn:0 {0}(1420,140)(1420,230){1}
wire w34;    //: /sn:0 {0}(790,317)(790,415)(1756,415){1}
wire w50;    //: /sn:0 {0}(1359,268)(1313,268){1}
wire w25;    //: /sn:0 {0}(-61,140)(-61,242){1}
wire w4;    //: /sn:0 {0}(1530,311)(1530,475)(1756,475){1}
wire w39;    //: /sn:0 {0}(883,193)(883,234){1}
wire w62;    //: /sn:0 {0}(806,140)(806,235){1}
wire w56;    //: /sn:0 {0}(1663,232)(1663,140){1}
wire w0;    //: /sn:0 {0}(556,140)(556,237){1}
wire w3;    //: /sn:0 {0}(495,275)(446,275){1}
wire w22;    //: /sn:0 {0}(648,193)(648,236){1}
wire w36;    //: /sn:0 {0}(293,321)(293,375)(1756,375){1}
wire w20;    //: /sn:0 {0}(55,140)(55,241){1}
wire w30;    //: /sn:0 {0}(-183,140)(-183,243){1}
wire w29;    //: /sn:0 {0}(907,316)(907,425)(1756,425){1}
wire w71;    //: /sn:0 {0}(1608,266)(1567,266){1}
wire w37;    //: /sn:0 {0}(409,320)(409,385)(1756,385){1}
wire w42;    //: /sn:0 {0}(827,272)(862,272){1}
wire w19;    //: /sn:0 {0}(1159,314)(1159,445)(1756,445){1}
wire w18;    //: /sn:0 {0}(120,278)(76,278){1}
wire w66;    //: /sn:0 {0}(1485,267)(1441,267){1}
wire w10;    //: /sn:0 {0}(425,140)(425,238){1}
wire w23;    //: /sn:0 {0}(-40,279)(-6,279){1}
wire w54;    //: /sn:0 {0}(1175,140)(1175,232){1}
wire w70;    //: /sn:0 {0}(1546,140)(1546,229){1}
wire w24;    //: /sn:0 {0}(1031,315)(1031,435)(1756,435){1}
wire w21;    //: /sn:0 {0}(15,193)(15,241){1}
wire w1;    //: /sn:0 {0}(516,193)(516,237){1}
wire w31;    //: /sn:0 {0}(-223,193)(-223,243){1}
wire w32;    //: /sn:0 {0}(-77,324)(-77,345)(1756,345){1}
wire w68;    //: /sn:0 {0}(672,318)(672,405)(1756,405){1}
wire w53;    //: /sn:0 {0}(1135,193)(1135,232){1}
wire w8;    //: /sn:0 {0}(248,277)(202,277){1}
wire w46;    //: /sn:0 {0}(1114,270)(1068,270){1}
wire w27;    //: /sn:0 {0}(1645,306)(1645,485)(1756,485){1}
wire w17;    //: /sn:0 {0}(688,236)(688,140){1}
wire w44;    //: /sn:0 {0}(1007,193)(1007,233){1}
wire w28;    //: /sn:0 {0}(-162,280)(-122,280){1}
wire w33;    //: /sn:0 {0}(39,323)(39,355)(1756,355){1}
wire w35;    //: /sn:0 {0}(165,322)(165,365)(1756,365){1}
wire w14;    //: /sn:0 {0}(1404,312)(1404,465)(1756,465){1}
wire w45;    //: /sn:0 {0}(1047,140)(1047,233){1}
wire w49;    //: /sn:0 {0}(1292,140)(1292,231){1}
wire w69;    //: /sn:0 {0}(1506,193)(1506,229){1}
wire w2;    //: /sn:0 {0}(627,274)(577,274){1}
wire w11;    //: /sn:0 {0}(385,193)(385,238){1}
wire w41;    //: /sn:0 {0}(986,271)(944,271){1}
wire w48;    //: /sn:0 {0}(1252,193)(1252,231){1}
wire w15;    //: /sn:0 {0}(181,140)(181,240){1}
wire w5;    //: /sn:0 {0}(309,140)(309,239){1}
wire w38;    //: /sn:0 {0}(540,319)(540,395)(1756,395){1}
wire w61;    //: /sn:0 {0}(766,193)(766,235){1}
wire w64;    //: /sn:0 {0}(1380,193)(1380,230){1}
wire w26;    //: /sn:0 {0}(-101,193)(-101,242){1}
wire w9;    //: /sn:0 {0}(1276,313)(1276,455)(1756,455){1}
wire w40;    //: /sn:0 {0}(923,140)(923,234){1}
wire w51;    //: /sn:0 {0}(1231,269)(1196,269){1}
wire w57;    //: /sn:0 {0}(1627,232)(1627,193){1}
//: enddecls

  FA g4 (.a(w21), .b(w20), .Cin(w18), .Cout(w23), .S(w33));   //: @(-5, 242) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  FA g8 (.a(w39), .b(w40), .Cin(w41), .Cout(w42), .S(w29));   //: @(863, 235) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  assign w69 = A[1]; //: TAP g44 @(1506,187) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  assign w16 = A[12]; //: TAP g16 @(141,187) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  FA g3 (.a(w16), .b(w15), .Cin(w8), .Cout(w18), .S(w35));   //: @(121, 241) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w40 = B[6]; //: TAP g47 @(923,134) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  assign w20 = B[13]; //: TAP g26 @(55,134) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  assign w6 = A[11]; //: TAP g17 @(269,187) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  FA g2 (.a(w11), .b(w10), .Cin(w3), .Cout(w7), .S(w37));   //: @(365, 239) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: comment g30 @(214,71) /sn:0
  //: /line:"Il Ripple Carry Adder (o RCA) è un modulo composto da tanti Full Adder collegati in serie, in base al numero di bit richiesti dall'operazione(in questo caso 8)."
  //: /end
  assign w10 = B[10]; //: TAP g23 @(425,134) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:1
  assign w5 = B[11]; //: TAP g24 @(309,134) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  FA g1 (.a(w6), .b(w5), .Cin(w7), .Cout(w8), .S(w36));   //: @(249, 240) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w39 = A[6]; //: TAP g39 @(883,187) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  assign S = {w13, w32, w33, w35, w36, w37, w38, w68, w34, w29, w24, w19, w9, w14, w4, w27}; //: CONCAT g29  @(1761,410) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  assign w65 = B[2]; //: TAP g51 @(1420,134) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  assign w11 = A[10]; //: TAP g18 @(385,187) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:1
  //: OUT g10 (S) @(1817,410) /sn:0 /w:[ 1 ]
  assign w15 = B[12]; //: TAP g25 @(181,134) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  assign w54 = B[4]; //: TAP g49 @(1175,134) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  FA g6 (.a(w31), .b(w30), .Cin(w28), .Cout(Cout), .S(w13));   //: @(-243, 244) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w49 = B[3]; //: TAP g50 @(1292,134) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  //: OUT g9 (Cout) @(1791,512) /sn:0 /w:[ 0 ]
  FA g35 (.a(w61), .b(w62), .Cin(w42), .Cout(w58), .S(w34));   //: @(746, 236) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  HA g7 (.a(w57), .b(w56), .Cout(w71), .S(w27));   //: @(1609, 233) /sz:(72, 72) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<0 ]
  assign w0 = B[9]; //: TAP g22 @(556,134) /sn:0 /R:1 /w:[ 0 20 19 ] /ss:1
  FA g31 (.a(w44), .b(w45), .Cin(w46), .Cout(w41), .S(w24));   //: @(987, 234) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g33 (.a(w53), .b(w54), .Cin(w51), .Cout(w46), .S(w19));   //: @(1115, 233) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g36 (.a(w64), .b(w65), .Cin(w66), .Cout(w50), .S(w14));   //: @(1360, 231) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w53 = A[4]; //: TAP g41 @(1135,187) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  assign w57 = A[0]; //: TAP g45 @(1627,187) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  assign w44 = A[5]; //: TAP g40 @(1007,187) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  assign w48 = A[3]; //: TAP g42 @(1252,187) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  assign w70 = B[1]; //: TAP g52 @(1546,134) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: IN g12 (B) @(-216,136) /sn:0 /w:[ 33 ]
  assign w30 = B[15]; //: TAP g28 @(-183,134) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:1
  FA g34 (.a(w22), .b(w17), .Cin(w58), .Cout(w2), .S(w68));   //: @(628, 237) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  assign w62 = B[7]; //: TAP g46 @(806,134) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  assign w26 = A[14]; //: TAP g14 @(-101,187) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:1
  //: IN g11 (A) @(-252,189) /sn:0 /w:[ 33 ]
  FA g5 (.a(w26), .b(w25), .Cin(w23), .Cout(w28), .S(w32));   //: @(-121, 243) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w17 = B[8]; //: TAP g21 @(688,134) /sn:0 /R:1 /w:[ 1 18 17 ] /ss:1
  assign w1 = A[9]; //: TAP g19 @(516,187) /sn:0 /R:1 /w:[ 0 20 19 ] /ss:1
  assign w22 = A[8]; //: TAP g20 @(648,187) /sn:0 /R:1 /w:[ 0 18 17 ] /ss:1
  FA g32 (.a(w48), .b(w49), .Cin(w50), .Cout(w51), .S(w9));   //: @(1232, 232) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w21 = A[13]; //: TAP g15 @(15,187) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  FA g0 (.a(w1), .b(w0), .Cin(w2), .Cout(w3), .S(w38));   //: @(496, 238) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w61 = A[7]; //: TAP g38 @(766,187) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  assign w64 = A[2]; //: TAP g43 @(1380,187) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  assign w25 = B[14]; //: TAP g27 @(-61,134) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:1
  assign w45 = B[5]; //: TAP g48 @(1047,134) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  FA g37 (.a(w69), .b(w70), .Cin(w71), .Cout(w66), .S(w4));   //: @(1486, 230) /sz:(80, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w31 = A[15]; //: TAP g13 @(-223,187) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:1
  assign w56 = B[0]; //: TAP g53 @(1663,134) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin NandEXOR
module NandEXOR(in2, out, in1);
//: interface  /sz:(99, 64) /bd:[ Li0>in2(44/64) Li1>in1(16/64) Ro0<out(27/64) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(280,341)(280,412){1}
//: {2}(278,414)(155,414)(155,643){3}
//: {4}(280,416)(280,430)(280,430)(280,451){5}
output out;    //: /sn:0 {0}(184,921)(184,971){1}
input in2;    //: /sn:0 {0}(109,341)(109,353)(109,353)(109,367){1}
//: {2}(111,369)(232,369)(232,643){3}
//: {4}(109,371)(109,451){5}
wire w13;    //: /sn:0 {0}(252,727)(252,788)(203,788)(203,837){1}
wire w7;    //: /sn:0 {0}(275,546)(275,590)(275,590)(275,643){1}
wire w12;    //: /sn:0 {0}(169,837)(169,785)(128,785)(128,732){1}
wire w9;    //: /sn:0 {0}(114,551)(114,643){1}
//: enddecls

  MyNAND g4 (.in1(w13), .in2(w12), .out(out));   //: @(151, 838) /sz:(70, 82) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 ]
  //: comment g8 @(70,-24) /sn:0
  //: /line:"La tabella di verità della porta EXOR è:"
  //: /line:""
  //: /line:" a | b | a(+)b"
  //: /line:"--------------"
  //: /line:" 0 | 0 |   0"
  //: /line:" 0 | 1 |   1"
  //: /line:" 1 | 0 |   1"
  //: /line:" 1 | 1 |   0"
  //: /line:""
  //: /line:"Traducibile in: a'b + ab'"
  //: /line:" "
  //: /line:" -> considerando a'b = x , ab' = y"
  //: /line:" -> De Morgan: x + y = (x' y')'"
  //: /line:" -> ((a'b)'(ab')')'"
  //: /end
  MyNAND g3 (.in1(in1), .in2(w9), .out(w12));   //: @(90, 644) /sz:(75, 87) /R:3 /sn:0 /p:[ Ti0>3 Ti1>1 Bo0<1 ]
  MyNAND g2 (.in1(w7), .in2(in2), .out(w13));   //: @(212, 644) /sz:(73, 82) /R:3 /sn:0 /p:[ Ti0>1 Ti1>3 Bo0<0 ]
  NandNOT g1 (.in1(in1), .out(w7));   //: @(243, 452) /sz:(52, 93) /R:3 /sn:0 /p:[ Ti0>5 Bo0<0 ]
  //: joint g10 (in1) @(280, 414) /w:[ -1 1 2 4 ]
  //: IN g6 (in2) @(109,339) /sn:0 /R:3 /w:[ 0 ]
  //: joint g9 (in2) @(109, 369) /w:[ 2 1 -1 4 ]
  //: OUT g7 (out) @(184,968) /sn:0 /R:3 /w:[ 1 ]
  //: IN g5 (in1) @(280,339) /sn:0 /R:3 /w:[ 0 ]
  NandNOT g0 (.in1(in2), .out(w9));   //: @(82, 452) /sz:(53, 98) /R:3 /sn:0 /p:[ Ti0>5 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin NandOR
module NandOR(in1, out, in2);
//: interface  /sz:(87, 64) /bd:[ Li0>in1(11/64) Li1>in2(48/64) Ro0<out(28/64) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(315,252)(315,208)(354,208){1}
//: {2}(356,206)(356,183){3}
//: {4}(356,210)(356,252){5}
output out;    //: /sn:0 {0}(264,530)(264,490){1}
input in2;    //: /sn:0 {0}(218,258)(218,215)(177,215){1}
//: {2}(175,217)(175,258){3}
//: {4}(175,213)(175,180){5}
wire w0;    //: /sn:0 {0}(312,341)(312,381)(289,381)(289,401){1}
wire w1;    //: /sn:0 {0}(242,401)(242,381)(218,381)(218,347){1}
//: enddecls

  //: IN g4 (in1) @(356,181) /sn:0 /R:3 /w:[ 3 ]
  //: OUT g8 (out) @(264,527) /sn:0 /R:3 /w:[ 0 ]
  MyNAND g3 (.in2(in1), .in1(in1), .out(w0));   //: @(299, 253) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>0 Ti1>5 Bo0<0 ]
  MyNAND g2 (.in2(in2), .in1(in2), .out(w1));   //: @(162, 259) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>3 Ti1>0 Bo0<1 ]
  MyNAND g1 (.in2(w1), .in1(w0), .out(out));   //: @(231, 402) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 ]
  //: IN g6 (in2) @(175,178) /sn:0 /R:3 /w:[ 5 ]
  //: joint g7 (in2) @(175, 215) /w:[ 2 1 4 -1 ]
  //: joint g5 (in1) @(356, 208) /w:[ -1 2 1 4 ]
  //: comment g0 @(134,-85) /sn:0
  //: /line:"L'OR è una porta logica elementare. "
  //: /line:"La sua tabella di verità è:"
  //: /line:""
  //: /line:" a | b | a+b"
  //: /line:" -----------"
  //: /line:" 0 | 0 | 0"
  //: /line:" 0 | 1 | 1"
  //: /line:" 1 | 0 | 1"
  //: /line:" 1 | 1 | 1"
  //: /line:""
  //: /line:"In logica NAND abbiamo: a+b -> ((aa)' (bb)')'"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin MyNAND
module MyNAND(out, in1, in2);
//: interface  /sz:(87, 64) /bd:[ Li0>in2(47/64) Li1>in1(16/64) Ro0<out(24/64) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(261,211)(302,211){1}
//: {2}(306,211)(322,211){3}
//: {4}(304,213)(304,290)(363,290){5}
supply1 w12;    //: /sn:0 {0}(375,158)(375,187){1}
//: {2}(377,189)(403,189)(403,204){3}
//: {4}(373,189)(336,189)(336,203){5}
supply0 w10;    //: /sn:0 {0}(377,383)(377,355){1}
output out;    //: /sn:0 {0}(377,282)(377,264){1}
//: {2}(379,262)(481,262){3}
//: {4}(377,260)(377,238){5}
//: {6}(379,236)(403,236)(403,221){7}
//: {8}(375,236)(336,236)(336,220){9}
input in2;    //: /sn:0 {0}(389,212)(345,212)(345,260){1}
//: {2}(343,262)(246,262){3}
//: {4}(345,264)(345,346)(363,346){5}
wire w6;    //: /sn:0 {0}(377,299)(377,338){1}
//: enddecls

  _GGNMOS #(2, 1) g4 (.Z(out), .S(w6), .G(in1));   //: @(371,290) /sn:0 /w:[ 0 0 5 ]
  //: joint g8 (w12) @(375, 189) /w:[ 2 1 4 -1 ]
  _GGNMOS #(2, 1) g3 (.Z(w6), .S(w10), .G(in2));   //: @(371,346) /sn:0 /w:[ 1 1 5 ]
  _GGPMOS #(2, 1) g2 (.Z(out), .S(w12), .G(in2));   //: @(397,212) /sn:0 /w:[ 7 3 0 ]
  _GGPMOS #(2, 1) g1 (.Z(out), .S(w12), .G(in1));   //: @(330,211) /sn:0 /w:[ 9 5 3 ]
  //: joint g10 (out) @(377, 262) /w:[ 2 4 -1 1 ]
  //: VDD g6 (w12) @(386,158) /sn:0 /w:[ 0 ]
  //: joint g7 (out) @(377, 236) /w:[ 6 -1 8 5 ]
  //: OUT g9 (out) @(478,262) /sn:0 /w:[ 3 ]
  //: joint g12 (in1) @(304, 211) /w:[ 2 -1 1 4 ]
  //: GROUND g5 (w10) @(377,389) /sn:0 /w:[ 0 ]
  //: IN g11 (in1) @(259,211) /sn:0 /w:[ 0 ]
  //: joint g14 (in2) @(345, 262) /w:[ -1 1 2 4 ]
  //: comment g0 @(185,-82) /sn:0
  //: /line:"Il Nand implementa un NOT AND."
  //: /line:"È una porta funzionalmente completa."
  //: /line:""
  //: /line:""
  //: /line:" A | B | AB | (AB)'"
  //: /line:"--------------------"
  //: /line:" 0 | 0 |  0 |  1"
  //: /line:" 0 | 1 |  0 |  1"
  //: /line:" 1 | 0 |  0 |  1"
  //: /line:" 1 | 1 |  1 |  0"
  //: /line:""
  //: /line:"Per il NOR è sufficiente invertire gli NMOS con i PMOS"
  //: /end
  //: IN g13 (in2) @(244,262) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX
module MUX(B, A, Cin, Y);
//: interface  /sz:(121, 48) /bd:[ Ti0>A(36/121) Ti1>B(86/121) Li0>Cin(24/48) Bo0<Y(63/121) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(551,16)(551,226){1}
input A;    //: /sn:0 {0}(352,11)(352,118)(352,118)(352,226){1}
input Cin;    //: /sn:0 {0}(379,78)(379,45)(403,45){1}
//: {2}(407,45)(515,45)(515,226){3}
//: {4}(405,43)(405,30)(405,30)(405,16){5}
//: {6}(405,47)(405,78){7}
output Y;    //: /sn:0 {0}(456,461)(456,523){1}
wire w8;    //: /sn:0 {0}(437,372)(437,333)(375,333)(375,315){1}
wire w2;    //: /sn:0 {0}(469,372)(469,332)(534,332)(534,316){1}
wire w5;    //: /sn:0 {0}(395,167)(395,196)(395,196)(395,226){1}
//: enddecls

  //: IN g4 (B) @(551,14) /sn:0 /R:3 /w:[ 0 ]
  //: IN g8 (A) @(352,9) /sn:0 /R:3 /w:[ 0 ]
  MyNAND g3 (.in2(w8), .in1(w2), .out(Y));   //: @(421, 373) /sz:(64, 87) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  MyNAND g2 (.in2(Cin), .in1(B), .out(w2));   //: @(497, 227) /sz:(69, 88) /R:3 /sn:0 /p:[ Ti0>3 Ti1>1 Bo0<1 ]
  MyNAND g1 (.in2(Cin), .in1(Cin), .out(w5));   //: @(361, 79) /sz:(61, 87) /R:3 /sn:0 /p:[ Ti0>0 Ti1>7 Bo0<0 ]
  //: IN g6 (Cin) @(405,14) /sn:0 /R:3 /w:[ 5 ]
  //: joint g9 (Cin) @(405, 45) /w:[ 2 4 1 6 ]
  //: OUT g5 (Y) @(456,520) /sn:0 /R:3 /w:[ 1 ]
  MyNAND g0 (.in2(A), .in1(w5), .out(w8));   //: @(336, 227) /sz:(71, 87) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin HS
module HS(D, B, Pr, A);
//: interface  /sz:(125, 46) /bd:[ Ti0>A(20/125) Ti1>B(90/125) Lo0<Pr(16/46) Bo0<D(20/125) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(335,174)(335,-1)(394,-1){1}
//: {2}(396,1)(396,174){3}
//: {4}(396,-3)(396,-39){5}
input A;    //: /sn:0 {0}(297,15)(297,-14)(435,-14){1}
//: {2}(437,-12)(437,174){3}
//: {4}(437,-16)(437,-39){5}
output Pr;    //: /sn:0 {0}(318,458)(318,438)(318,438)(318,416){1}
output D;    //: /sn:0 {0}(417,275)(417,458){1}
wire w1;    //: /sn:0 {0}(300,110)(300,174){1}
wire w5;    //: /sn:0 {0}(318,277)(318,321){1}
//: enddecls

  MyNAND g4 (.in2(w1), .in1(B), .out(w5));   //: @(281, 175) /sz:(64, 101) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 ]
  //: OUT g8 (D) @(417,455) /sn:0 /R:3 /w:[ 1 ]
  NandNOT g3 (.in1(A), .out(w1));   //: @(263, 16) /sz:(48, 93) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  NandEXOR g2 (.in2(B), .in1(A), .out(D));   //: @(380, 175) /sz:(64, 99) /R:3 /sn:0 /p:[ Ti0>3 Ti1>3 Bo0<0 ]
  //: IN g1 (B) @(396,-41) /sn:0 /R:3 /w:[ 5 ]
  //: joint g6 (A) @(437, -14) /w:[ 2 -1 4 1 ]
  //: joint g7 (B) @(396, -1) /w:[ 2 -1 4 1 ]
  //: OUT g9 (Pr) @(318,455) /sn:0 /R:3 /w:[ 0 ]
  NandNOT g5 (.in1(w5), .out(Pr));   //: @(286, 322) /sz:(48, 93) /R:3 /sn:0 /p:[ Ti0>1 Bo0<1 ]
  //: IN g0 (A) @(437,-41) /sn:0 /R:3 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(b, a, Cout, S, Cin);
//: interface  /sz:(82, 75) /bd:[ Ti0>a(29/82) Ti1>b(57/82) Ri0>Cin(37/75) Lo0<Cout(38/75) Bo0<S(41/82) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(253,228)(253,258){1}
input Cin;    //: /sn:0 {0}(283,398)(283,228){1}
output Cout;    //: /sn:0 {0}(162,571)(162,551)(162,551)(162,533){1}
input a;    //: /sn:0 {0}(221,228)(221,258){1}
output S;    //: /sn:0 {0}(270,571)(270,474){1}
wire w4;    //: /sn:0 {0}(227,432)(179,432)(179,447){1}
wire w3;    //: /sn:0 {0}(255,398)(255,364)(229,364)(229,332){1}
wire w2;    //: /sn:0 {0}(193,292)(146,292)(146,447){1}
//: enddecls

  //: IN g4 (b) @(253,226) /sn:0 /R:3 /w:[ 0 ]
  NandOR g8 (.in1(w4), .in2(w2), .out(Cout));   //: @(130, 448) /sz:(64, 84) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  //: IN g3 (a) @(221,226) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g2 (Cout) @(162,568) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g1 (S) @(270,568) /sn:0 /R:3 /w:[ 0 ]
  HA g6 (.a(a), .b(b), .Cout(w2), .S(w3));   //: @(194, 259) /sz:(81, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<1 ]
  HA g7 (.a(w3), .b(Cin), .Cout(w4), .S(S));   //: @(229, 399) /sz:(89, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  //: IN g5 (Cin) @(283,226) /sn:0 /R:3 /w:[ 1 ]
  //: comment g0 @(-46,-40) /sn:0
  //: /line:"Il FULL ADDER (FA) permette di eseguire una somma tra singoli bit, di prendere in ingresso ed ventualmente propagare il riporto."
  //: /line:""
  //: /line:"La sua tabella della verità è:"
  //: /line:""
  //: /line:" a | b | Cin | S | Cout"
  //: /line:"------------------------"
  //: /line:" 0 | 0 |  0  | 0 |  0"
  //: /line:" 0 | 0 |  1  | 1 |  0"
  //: /line:" 0 | 1 |  0  | 1 |  0"
  //: /line:" 0 | 1 |  1  | 0 |  1"
  //: /line:" 1 | 0 |  0  | 1 |  0"
  //: /line:" 1 | 0 |  1  | 0 |  1"
  //: /line:" 1 | 1 |  0  | 0 |  1"
  //: /line:" 1 | 1 |  1  | 1 |  1"
  //: /end

endmodule
//: /netlistEnd

